module multiplier( input [127:0] x , output [127:0] y );
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 ,
    n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 ,
    n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 ,
    n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 ,
    n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 ,
    n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 ,
    n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 ,
    n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 ,
    n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 ,
    n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 ,
    n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 ,
    n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 ,
    n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 ,
    n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 ,
    n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 ,
    n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 ,
    n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 ,
    n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 ,
    n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 ,
    n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 ,
    n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 ,
    n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 ,
    n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 ,
    n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 ,
    n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 ,
    n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 ,
    n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 ,
    n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 ,
    n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 ,
    n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 ,
    n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 ,
    n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 ,
    n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 ,
    n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 ,
    n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 ;
  assign n129 = x[0] & x[64] ;
  assign n27784 = ~n129 ;
  assign n22786 = x[2] & n27784 ;
  assign n258 = x[64] & x[65] ;
  assign n6436 = x[64] | x[65] ;
  assign n27785 = ~n258 ;
  assign n6437 = n27785 & n6436 ;
  assign n278 = x[1] & x[2] ;
  assign n19653 = x[1] | x[2] ;
  assign n27786 = ~n278 ;
  assign n19654 = n27786 & n19653 ;
  assign n19656 = x[0] & n19654 ;
  assign n19658 = n6437 & n19656 ;
  assign n27787 = ~x[0] ;
  assign n19829 = n27787 & x[1] ;
  assign n22787 = x[64] & n19829 ;
  assign n27788 = ~n19654 ;
  assign n19655 = x[0] & n27788 ;
  assign n22788 = x[65] & n19655 ;
  assign n22789 = n22787 | n22788 ;
  assign n22790 = n19658 | n22789 ;
  assign n27789 = ~n22790 ;
  assign n22791 = x[2] & n27789 ;
  assign n27790 = ~x[2] ;
  assign n22792 = n27790 & n22790 ;
  assign n22793 = n22791 | n22792 ;
  assign n22794 = n22786 | n22793 ;
  assign n22795 = n22786 & n22793 ;
  assign n27791 = ~n22795 ;
  assign n130 = n22794 & n27791 ;
  assign n27792 = ~x[66] ;
  assign n6461 = x[64] & n27792 ;
  assign n6462 = x[65] & n6461 ;
  assign n259 = x[65] & x[66] ;
  assign n6463 = x[65] | x[66] ;
  assign n27793 = ~n259 ;
  assign n6464 = n27793 & n6463 ;
  assign n6465 = n258 | n6464 ;
  assign n27794 = ~n6462 ;
  assign n6466 = n27794 & n6465 ;
  assign n19683 = n6466 & n19656 ;
  assign n19722 = n27787 & n19654 ;
  assign n27795 = ~x[1] ;
  assign n19723 = n27795 & n19722 ;
  assign n19765 = x[64] & n19723 ;
  assign n19850 = x[65] & n19829 ;
  assign n22796 = n19765 | n19850 ;
  assign n22797 = x[66] & n19655 ;
  assign n22798 = n22796 | n22797 ;
  assign n22799 = n19683 | n22798 ;
  assign n27796 = ~n22799 ;
  assign n22800 = x[2] & n27796 ;
  assign n22801 = n27790 & n22799 ;
  assign n22802 = n22800 | n22801 ;
  assign n22803 = n22795 | n22802 ;
  assign n22804 = n22795 & n22802 ;
  assign n27797 = ~n22804 ;
  assign n131 = n22803 & n27797 ;
  assign n276 = x[2] & x[3] ;
  assign n18323 = x[2] | x[3] ;
  assign n27798 = ~n276 ;
  assign n18324 = n27798 & n18323 ;
  assign n21799 = x[64] & n18324 ;
  assign n453 = x[64] | x[66] ;
  assign n454 = x[65] & n453 ;
  assign n27653 = x[66] & x[67] ;
  assign n455 = x[66] | x[67] ;
  assign n27799 = ~n27653 ;
  assign n456 = n27799 & n455 ;
  assign n457 = n454 | n456 ;
  assign n458 = n454 & n456 ;
  assign n27800 = ~n458 ;
  assign n6494 = n457 & n27800 ;
  assign n19709 = n6494 & n19656 ;
  assign n19724 = x[65] & n19723 ;
  assign n19836 = x[66] & n19829 ;
  assign n22777 = n19724 | n19836 ;
  assign n22778 = x[67] & n19655 ;
  assign n22779 = n22777 | n22778 ;
  assign n22780 = n19709 | n22779 ;
  assign n27801 = ~n22780 ;
  assign n22781 = x[2] & n27801 ;
  assign n22782 = n27790 & n22780 ;
  assign n22783 = n22781 | n22782 ;
  assign n27802 = ~n22783 ;
  assign n22784 = n21799 & n27802 ;
  assign n27803 = ~n21799 ;
  assign n22805 = n27803 & n22783 ;
  assign n22806 = n22784 | n22805 ;
  assign n22807 = n22804 & n22806 ;
  assign n27621 = n22804 | n22806 ;
  assign n27804 = ~n22807 ;
  assign n132 = n27804 & n27621 ;
  assign n459 = n27653 | n458 ;
  assign n27145 = x[67] & x[68] ;
  assign n460 = x[67] | x[68] ;
  assign n27805 = ~n27145 ;
  assign n461 = n27805 & n460 ;
  assign n462 = n459 & n461 ;
  assign n6407 = n459 | n461 ;
  assign n27806 = ~n462 ;
  assign n6408 = n27806 & n6407 ;
  assign n19693 = n6408 & n19656 ;
  assign n19735 = x[66] & n19723 ;
  assign n19874 = x[67] & n19829 ;
  assign n22766 = n19735 | n19874 ;
  assign n22767 = x[68] & n19655 ;
  assign n22768 = n22766 | n22767 ;
  assign n22769 = n19693 | n22768 ;
  assign n22770 = x[2] | n22769 ;
  assign n22771 = x[2] & n22769 ;
  assign n27807 = ~n22771 ;
  assign n22772 = n22770 & n27807 ;
  assign n21800 = x[5] & n27803 ;
  assign n277 = x[4] & x[5] ;
  assign n18325 = x[4] | x[5] ;
  assign n27808 = ~n277 ;
  assign n18326 = n27808 & n18325 ;
  assign n18392 = n18324 & n18326 ;
  assign n18400 = n6437 & n18392 ;
  assign n275 = x[3] & x[4] ;
  assign n18321 = x[3] | x[4] ;
  assign n27809 = ~n275 ;
  assign n18322 = n27809 & n18321 ;
  assign n27810 = ~n18324 ;
  assign n18514 = n18322 & n27810 ;
  assign n21801 = x[64] & n18514 ;
  assign n27811 = ~n18326 ;
  assign n18327 = n18324 & n27811 ;
  assign n21802 = x[65] & n18327 ;
  assign n21803 = n21801 | n21802 ;
  assign n21804 = n18400 | n21803 ;
  assign n27812 = ~n21804 ;
  assign n21805 = x[5] & n27812 ;
  assign n27813 = ~x[5] ;
  assign n21806 = n27813 & n21804 ;
  assign n21807 = n21805 | n21806 ;
  assign n21808 = n21800 | n21807 ;
  assign n21809 = n21800 & n21807 ;
  assign n27814 = ~n21809 ;
  assign n22773 = n21808 & n27814 ;
  assign n22774 = n22772 & n22773 ;
  assign n22775 = n22772 | n22773 ;
  assign n27815 = ~n22774 ;
  assign n22776 = n27815 & n22775 ;
  assign n22785 = n21799 & n22783 ;
  assign n22808 = n22785 | n22807 ;
  assign n22809 = n22776 & n22808 ;
  assign n27623 = n22776 | n22808 ;
  assign n27816 = ~n22809 ;
  assign n133 = n27816 & n27623 ;
  assign n463 = n27145 | n462 ;
  assign n27652 = x[68] & x[69] ;
  assign n464 = x[68] | x[69] ;
  assign n27817 = ~n27652 ;
  assign n465 = n27817 & n464 ;
  assign n466 = n463 | n465 ;
  assign n467 = n463 & n465 ;
  assign n27818 = ~n467 ;
  assign n6379 = n466 & n27818 ;
  assign n19667 = n6379 & n19656 ;
  assign n19725 = x[67] & n19723 ;
  assign n19882 = x[68] & n19829 ;
  assign n22754 = n19725 | n19882 ;
  assign n22755 = x[69] & n19655 ;
  assign n22756 = n22754 | n22755 ;
  assign n22757 = n19667 | n22756 ;
  assign n27819 = ~n22757 ;
  assign n22758 = x[2] & n27819 ;
  assign n22759 = n27790 & n22757 ;
  assign n22760 = n22758 | n22759 ;
  assign n18455 = n6466 & n18392 ;
  assign n21810 = x[66] & n18327 ;
  assign n18328 = n27810 & n18326 ;
  assign n27820 = ~n18322 ;
  assign n18329 = n27820 & n18328 ;
  assign n21811 = x[64] & n18329 ;
  assign n21812 = x[65] & n18514 ;
  assign n21813 = n21811 | n21812 ;
  assign n21814 = n21810 | n21813 ;
  assign n21815 = n18455 | n21814 ;
  assign n27821 = ~n21815 ;
  assign n21816 = x[5] & n27821 ;
  assign n21817 = n27813 & n21815 ;
  assign n21818 = n21816 | n21817 ;
  assign n21819 = n21809 | n21818 ;
  assign n21820 = n21809 & n21818 ;
  assign n27822 = ~n21820 ;
  assign n22761 = n21819 & n27822 ;
  assign n27823 = ~n22760 ;
  assign n22762 = n27823 & n22761 ;
  assign n27824 = ~n22761 ;
  assign n22764 = n22760 & n27824 ;
  assign n22765 = n22762 | n22764 ;
  assign n22810 = n22774 | n22809 ;
  assign n22811 = n22765 | n22810 ;
  assign n22812 = n22765 & n22810 ;
  assign n27825 = ~n22812 ;
  assign n134 = n22811 & n27825 ;
  assign n22763 = n22760 & n22761 ;
  assign n22813 = n22763 | n22812 ;
  assign n273 = x[5] & x[6] ;
  assign n15240 = x[5] | x[6] ;
  assign n27826 = ~n273 ;
  assign n15241 = n27826 & n15240 ;
  assign n20716 = x[64] & n15241 ;
  assign n27827 = ~n20716 ;
  assign n21822 = n27827 & n21820 ;
  assign n22145 = n20716 & n27822 ;
  assign n22146 = n21822 | n22145 ;
  assign n18456 = n6494 & n18392 ;
  assign n18355 = x[65] & n18329 ;
  assign n18574 = x[66] & n18514 ;
  assign n21825 = n18355 | n18574 ;
  assign n21826 = x[67] & n18327 ;
  assign n21827 = n21825 | n21826 ;
  assign n21828 = n18456 | n21827 ;
  assign n27828 = ~n21828 ;
  assign n21830 = x[5] & n27828 ;
  assign n22147 = n27813 & n21828 ;
  assign n22148 = n21830 | n22147 ;
  assign n22149 = n22146 | n22148 ;
  assign n22150 = n22146 & n22148 ;
  assign n27829 = ~n22150 ;
  assign n22744 = n22149 & n27829 ;
  assign n468 = n27652 | n467 ;
  assign n27074 = x[69] & x[70] ;
  assign n469 = x[69] | x[70] ;
  assign n27830 = ~n27074 ;
  assign n5973 = n27830 & n469 ;
  assign n5974 = n468 & n5973 ;
  assign n5975 = n468 | n5973 ;
  assign n27831 = ~n5974 ;
  assign n5976 = n27831 & n5975 ;
  assign n19702 = n5976 & n19656 ;
  assign n19784 = x[68] & n19723 ;
  assign n19834 = x[69] & n19829 ;
  assign n22745 = n19784 | n19834 ;
  assign n22746 = x[70] & n19655 ;
  assign n22747 = n22745 | n22746 ;
  assign n22748 = n19702 | n22747 ;
  assign n27832 = ~n22748 ;
  assign n22749 = x[2] & n27832 ;
  assign n22750 = n27790 & n22748 ;
  assign n22751 = n22749 | n22750 ;
  assign n27833 = ~n22751 ;
  assign n22752 = n22744 & n27833 ;
  assign n27834 = ~n22744 ;
  assign n22814 = n27834 & n22751 ;
  assign n22815 = n22752 | n22814 ;
  assign n22816 = n22813 & n22815 ;
  assign n27626 = n22813 | n22815 ;
  assign n27835 = ~n22816 ;
  assign n135 = n27835 & n27626 ;
  assign n22753 = n22744 & n22751 ;
  assign n22817 = n22753 | n22816 ;
  assign n470 = n468 & n469 ;
  assign n471 = n27074 | n470 ;
  assign n27655 = x[70] & x[71] ;
  assign n472 = x[70] | x[71] ;
  assign n27836 = ~n27655 ;
  assign n473 = n27836 & n472 ;
  assign n474 = n471 | n473 ;
  assign n475 = n471 & n473 ;
  assign n27837 = ~n475 ;
  assign n4790 = n474 & n27837 ;
  assign n19660 = n4790 & n19656 ;
  assign n19727 = x[69] & n19723 ;
  assign n19842 = x[70] & n19829 ;
  assign n22734 = n19727 | n19842 ;
  assign n22735 = x[71] & n19655 ;
  assign n22736 = n22734 | n22735 ;
  assign n22737 = n19660 | n22736 ;
  assign n27838 = ~n22737 ;
  assign n22738 = x[2] & n27838 ;
  assign n22739 = n27790 & n22737 ;
  assign n22740 = n22738 | n22739 ;
  assign n18423 = n6408 & n18392 ;
  assign n18371 = x[66] & n18329 ;
  assign n18563 = x[67] & n18514 ;
  assign n21786 = n18371 | n18563 ;
  assign n21787 = x[68] & n18327 ;
  assign n21788 = n21786 | n21787 ;
  assign n21789 = n18423 | n21788 ;
  assign n27839 = ~n21789 ;
  assign n21790 = x[5] & n27839 ;
  assign n21792 = n27813 & n21789 ;
  assign n21793 = n21790 | n21792 ;
  assign n20717 = x[8] & n27827 ;
  assign n274 = x[7] & x[8] ;
  assign n15242 = x[7] | x[8] ;
  assign n27840 = ~n274 ;
  assign n15243 = n27840 & n15242 ;
  assign n15308 = n15241 & n15243 ;
  assign n15369 = n6437 & n15308 ;
  assign n272 = x[6] & x[7] ;
  assign n15238 = x[6] | x[7] ;
  assign n27841 = ~n272 ;
  assign n15239 = n27841 & n15238 ;
  assign n27842 = ~n15241 ;
  assign n16288 = n15239 & n27842 ;
  assign n20718 = x[64] & n16288 ;
  assign n27843 = ~n15243 ;
  assign n15244 = n15241 & n27843 ;
  assign n20719 = x[65] & n15244 ;
  assign n20720 = n20718 | n20719 ;
  assign n20721 = n15369 | n20720 ;
  assign n27844 = ~n20721 ;
  assign n20722 = x[8] & n27844 ;
  assign n27845 = ~x[8] ;
  assign n20723 = n27845 & n20721 ;
  assign n20724 = n20722 | n20723 ;
  assign n20725 = n20717 | n20724 ;
  assign n20726 = n20717 & n20724 ;
  assign n27846 = ~n20726 ;
  assign n21794 = n20725 & n27846 ;
  assign n27847 = ~n21793 ;
  assign n21795 = n27847 & n21794 ;
  assign n27848 = ~n21794 ;
  assign n21797 = n21793 & n27848 ;
  assign n21798 = n21795 | n21797 ;
  assign n21821 = n20716 & n21820 ;
  assign n21823 = n20716 | n21820 ;
  assign n27849 = ~n21821 ;
  assign n21824 = n27849 & n21823 ;
  assign n21829 = x[5] | n21828 ;
  assign n21831 = x[5] & n21828 ;
  assign n27850 = ~n21831 ;
  assign n21832 = n21829 & n27850 ;
  assign n21833 = n21824 & n21832 ;
  assign n21834 = n21821 | n21833 ;
  assign n21835 = n21798 | n21834 ;
  assign n21836 = n21798 & n21834 ;
  assign n27851 = ~n21836 ;
  assign n22741 = n21835 & n27851 ;
  assign n27852 = ~n22740 ;
  assign n22742 = n27852 & n22741 ;
  assign n27853 = ~n22741 ;
  assign n22818 = n22740 & n27853 ;
  assign n22819 = n22742 | n22818 ;
  assign n22820 = n22817 | n22819 ;
  assign n22821 = n22817 & n22819 ;
  assign n27854 = ~n22821 ;
  assign n136 = n22820 & n27854 ;
  assign n15370 = n6466 & n15308 ;
  assign n15245 = n27842 & n15243 ;
  assign n27855 = ~n15239 ;
  assign n15246 = n27855 & n15245 ;
  assign n15285 = x[64] & n15246 ;
  assign n17274 = x[65] & n16288 ;
  assign n20727 = n15285 | n17274 ;
  assign n20728 = x[66] & n15244 ;
  assign n20729 = n20727 | n20728 ;
  assign n20730 = n15370 | n20729 ;
  assign n27856 = ~n20730 ;
  assign n20731 = x[8] & n27856 ;
  assign n20732 = n27845 & n20730 ;
  assign n20733 = n20731 | n20732 ;
  assign n20734 = n20726 & n20733 ;
  assign n20748 = n20726 | n20733 ;
  assign n27857 = ~n20734 ;
  assign n21774 = n27857 & n20748 ;
  assign n18454 = n6379 & n18392 ;
  assign n18330 = x[67] & n18329 ;
  assign n18515 = x[68] & n18514 ;
  assign n21775 = n18330 | n18515 ;
  assign n21776 = x[69] & n18327 ;
  assign n21777 = n21775 | n21776 ;
  assign n21778 = n18454 | n21777 ;
  assign n27858 = ~n21778 ;
  assign n21779 = x[5] & n27858 ;
  assign n21780 = n27813 & n21778 ;
  assign n21781 = n21779 | n21780 ;
  assign n27859 = ~n21781 ;
  assign n21782 = n21774 & n27859 ;
  assign n27860 = ~n21774 ;
  assign n21784 = n27860 & n21781 ;
  assign n21785 = n21782 | n21784 ;
  assign n21791 = x[5] | n21789 ;
  assign n22140 = x[5] & n21789 ;
  assign n27861 = ~n22140 ;
  assign n22141 = n21791 & n27861 ;
  assign n22142 = n21794 & n22141 ;
  assign n22143 = n21794 | n22141 ;
  assign n27862 = ~n22142 ;
  assign n22144 = n27862 & n22143 ;
  assign n22151 = n21821 | n22150 ;
  assign n22152 = n22144 & n22151 ;
  assign n22153 = n22142 | n22152 ;
  assign n22154 = n21785 | n22153 ;
  assign n22155 = n21785 & n22153 ;
  assign n27863 = ~n22155 ;
  assign n22722 = n22154 & n27863 ;
  assign n476 = n27655 | n475 ;
  assign n27656 = x[71] & x[72] ;
  assign n477 = x[71] | x[72] ;
  assign n27864 = ~n27656 ;
  assign n478 = n27864 & n477 ;
  assign n27865 = ~n476 ;
  assign n479 = n27865 & n478 ;
  assign n27866 = ~n478 ;
  assign n3700 = n476 & n27866 ;
  assign n3701 = n479 | n3700 ;
  assign n19690 = n3701 & n19656 ;
  assign n19749 = x[70] & n19723 ;
  assign n19835 = x[71] & n19829 ;
  assign n22723 = n19749 | n19835 ;
  assign n22724 = x[72] & n19655 ;
  assign n22725 = n22723 | n22724 ;
  assign n22726 = n19690 | n22725 ;
  assign n27867 = ~n22726 ;
  assign n22727 = x[2] & n27867 ;
  assign n22728 = n27790 & n22726 ;
  assign n22729 = n22727 | n22728 ;
  assign n27868 = ~n22729 ;
  assign n22730 = n22722 & n27868 ;
  assign n27869 = ~n22722 ;
  assign n22732 = n27869 & n22729 ;
  assign n22733 = n22730 | n22732 ;
  assign n22743 = n22740 & n22741 ;
  assign n22822 = n22743 | n22821 ;
  assign n22823 = n22733 & n22822 ;
  assign n27629 = n22733 | n22822 ;
  assign n27870 = ~n22823 ;
  assign n137 = n27870 & n27629 ;
  assign n18393 = n5976 & n18392 ;
  assign n18376 = x[68] & n18329 ;
  assign n18520 = x[69] & n18514 ;
  assign n21759 = n18376 | n18520 ;
  assign n21760 = x[70] & n18327 ;
  assign n21761 = n21759 | n21760 ;
  assign n21762 = n18393 | n21761 ;
  assign n27871 = ~n21762 ;
  assign n21763 = x[5] & n27871 ;
  assign n21764 = n27813 & n21762 ;
  assign n21765 = n21763 | n21764 ;
  assign n15371 = n6494 & n15308 ;
  assign n15307 = x[65] & n15246 ;
  assign n17295 = x[66] & n16288 ;
  assign n20739 = n15307 | n17295 ;
  assign n20740 = x[67] & n15244 ;
  assign n20741 = n20739 | n20740 ;
  assign n20742 = n15371 | n20741 ;
  assign n27872 = ~n20742 ;
  assign n20743 = x[8] & n27872 ;
  assign n20744 = n27845 & n20742 ;
  assign n20745 = n20743 | n20744 ;
  assign n270 = x[8] & x[9] ;
  assign n12627 = x[8] | x[9] ;
  assign n27873 = ~n270 ;
  assign n12628 = n27873 & n12627 ;
  assign n19365 = x[64] & n12628 ;
  assign n27874 = ~n19365 ;
  assign n20736 = n27874 & n20734 ;
  assign n21154 = n19365 & n27857 ;
  assign n21155 = n20736 | n21154 ;
  assign n21156 = n20745 | n21155 ;
  assign n21157 = n20745 & n21155 ;
  assign n27875 = ~n21157 ;
  assign n21769 = n21156 & n27875 ;
  assign n27876 = ~n21765 ;
  assign n21770 = n27876 & n21769 ;
  assign n27877 = ~n21769 ;
  assign n21772 = n21765 & n27877 ;
  assign n21773 = n21770 | n21772 ;
  assign n21783 = n21774 & n21781 ;
  assign n21796 = n21793 & n21794 ;
  assign n21837 = n21796 | n21836 ;
  assign n21838 = n21785 & n21837 ;
  assign n21839 = n21783 | n21838 ;
  assign n21840 = n21773 | n21839 ;
  assign n21841 = n21773 & n21839 ;
  assign n27878 = ~n21841 ;
  assign n22710 = n21840 & n27878 ;
  assign n480 = n476 & n478 ;
  assign n481 = n27656 | n480 ;
  assign n27650 = x[72] & x[73] ;
  assign n482 = x[72] | x[73] ;
  assign n27879 = ~n27650 ;
  assign n3730 = n27879 & n482 ;
  assign n3731 = n481 | n3730 ;
  assign n3732 = n481 & n3730 ;
  assign n27880 = ~n3732 ;
  assign n3733 = n3731 & n27880 ;
  assign n19662 = n3733 & n19656 ;
  assign n19750 = x[71] & n19723 ;
  assign n19839 = x[72] & n19829 ;
  assign n22711 = n19750 | n19839 ;
  assign n22712 = x[73] & n19655 ;
  assign n22713 = n22711 | n22712 ;
  assign n22714 = n19662 | n22713 ;
  assign n27881 = ~n22714 ;
  assign n22715 = x[2] & n27881 ;
  assign n22716 = n27790 & n22714 ;
  assign n22717 = n22715 | n22716 ;
  assign n27882 = ~n22717 ;
  assign n22718 = n22710 & n27882 ;
  assign n27883 = ~n22710 ;
  assign n22720 = n27883 & n22717 ;
  assign n22721 = n22718 | n22720 ;
  assign n22731 = n22722 & n22729 ;
  assign n22824 = n22731 | n22823 ;
  assign n22825 = n22721 | n22824 ;
  assign n22826 = n22721 & n22824 ;
  assign n27884 = ~n22826 ;
  assign n138 = n22825 & n27884 ;
  assign n22719 = n22710 & n22717 ;
  assign n22827 = n22719 | n22826 ;
  assign n18448 = n4790 & n18392 ;
  assign n18370 = x[69] & n18329 ;
  assign n18552 = x[70] & n18514 ;
  assign n21746 = n18370 | n18552 ;
  assign n21747 = x[71] & n18327 ;
  assign n21748 = n21746 | n21747 ;
  assign n21749 = n18448 | n21748 ;
  assign n27885 = ~n21749 ;
  assign n21750 = x[5] & n27885 ;
  assign n21751 = n27813 & n21749 ;
  assign n21752 = n21750 | n21751 ;
  assign n20735 = n19365 & n20734 ;
  assign n21158 = n20735 | n21157 ;
  assign n15356 = n6408 & n15308 ;
  assign n15306 = x[66] & n15246 ;
  assign n17324 = x[67] & n16288 ;
  assign n20707 = n15306 | n17324 ;
  assign n20708 = x[68] & n15244 ;
  assign n20709 = n20707 | n20708 ;
  assign n20710 = n15356 | n20709 ;
  assign n27886 = ~n20710 ;
  assign n20711 = x[8] & n27886 ;
  assign n20712 = n27845 & n20710 ;
  assign n20713 = n20711 | n20712 ;
  assign n19366 = x[11] & n27874 ;
  assign n271 = x[10] & x[11] ;
  assign n12629 = x[10] | x[11] ;
  assign n27887 = ~n271 ;
  assign n12630 = n27887 & n12629 ;
  assign n12695 = n12628 & n12630 ;
  assign n12750 = n6437 & n12695 ;
  assign n269 = x[9] & x[10] ;
  assign n12625 = x[9] | x[10] ;
  assign n27888 = ~n269 ;
  assign n12626 = n27888 & n12625 ;
  assign n27889 = ~n12628 ;
  assign n13533 = n12626 & n27889 ;
  assign n19367 = x[64] & n13533 ;
  assign n27890 = ~n12630 ;
  assign n12631 = n12628 & n27890 ;
  assign n19368 = x[65] & n12631 ;
  assign n19369 = n19367 | n19368 ;
  assign n19370 = n12750 | n19369 ;
  assign n27891 = ~n19370 ;
  assign n19371 = x[11] & n27891 ;
  assign n27892 = ~x[11] ;
  assign n19372 = n27892 & n19370 ;
  assign n19373 = n19371 | n19372 ;
  assign n19374 = n19366 | n19373 ;
  assign n19375 = n19366 & n19373 ;
  assign n27893 = ~n19375 ;
  assign n20714 = n19374 & n27893 ;
  assign n20715 = n20713 & n20714 ;
  assign n20750 = n20713 | n20714 ;
  assign n27894 = ~n20715 ;
  assign n21159 = n27894 & n20750 ;
  assign n21160 = n21158 & n21159 ;
  assign n21753 = n21158 | n21159 ;
  assign n27895 = ~n21160 ;
  assign n21754 = n27895 & n21753 ;
  assign n21755 = n21752 & n21754 ;
  assign n21757 = n21752 | n21754 ;
  assign n27896 = ~n21755 ;
  assign n21758 = n27896 & n21757 ;
  assign n20737 = n19365 | n20734 ;
  assign n27897 = ~n20735 ;
  assign n20738 = n27897 & n20737 ;
  assign n27898 = ~n20745 ;
  assign n20747 = n20738 & n27898 ;
  assign n27899 = ~n20738 ;
  assign n21766 = n27899 & n20745 ;
  assign n21767 = n20747 | n21766 ;
  assign n21768 = n21765 & n21767 ;
  assign n21771 = n21765 & n21769 ;
  assign n22138 = n21765 | n21769 ;
  assign n27900 = ~n21771 ;
  assign n22139 = n27900 & n22138 ;
  assign n22156 = n21783 | n22155 ;
  assign n22157 = n22139 & n22156 ;
  assign n22158 = n21768 | n22157 ;
  assign n27901 = ~n22158 ;
  assign n22159 = n21758 & n27901 ;
  assign n27902 = ~n21758 ;
  assign n22699 = n27902 & n22158 ;
  assign n22700 = n22159 | n22699 ;
  assign n483 = n481 & n482 ;
  assign n484 = n27650 | n483 ;
  assign n26995 = x[73] & x[74] ;
  assign n485 = x[73] | x[74] ;
  assign n27903 = ~n26995 ;
  assign n2719 = n27903 & n485 ;
  assign n2720 = n484 & n2719 ;
  assign n2721 = n484 | n2719 ;
  assign n27904 = ~n2720 ;
  assign n2722 = n27904 & n2721 ;
  assign n19679 = n2722 & n19656 ;
  assign n19739 = x[72] & n19723 ;
  assign n19853 = x[73] & n19829 ;
  assign n22701 = n19739 | n19853 ;
  assign n22702 = x[74] & n19655 ;
  assign n22703 = n22701 | n22702 ;
  assign n22704 = n19679 | n22703 ;
  assign n27905 = ~n22704 ;
  assign n22705 = x[2] & n27905 ;
  assign n22706 = n27790 & n22704 ;
  assign n22707 = n22705 | n22706 ;
  assign n22708 = n22700 | n22707 ;
  assign n22709 = n22700 & n22707 ;
  assign n27906 = ~n22709 ;
  assign n22828 = n22708 & n27906 ;
  assign n22829 = n22827 & n22828 ;
  assign n27632 = n22827 | n22828 ;
  assign n27907 = ~n22829 ;
  assign n139 = n27907 & n27632 ;
  assign n22830 = n22709 | n22829 ;
  assign n18394 = n3701 & n18392 ;
  assign n18334 = x[70] & n18329 ;
  assign n18517 = x[71] & n18514 ;
  assign n21737 = n18334 | n18517 ;
  assign n21738 = x[72] & n18327 ;
  assign n21739 = n21737 | n21738 ;
  assign n21740 = n18394 | n21739 ;
  assign n27908 = ~n21740 ;
  assign n21741 = x[5] & n27908 ;
  assign n21742 = n27813 & n21740 ;
  assign n21743 = n21741 | n21742 ;
  assign n12700 = n6466 & n12695 ;
  assign n12632 = n27889 & n12630 ;
  assign n27909 = ~n12626 ;
  assign n12633 = n27909 & n12632 ;
  assign n12693 = x[64] & n12633 ;
  assign n14383 = x[65] & n13533 ;
  assign n19376 = n12693 | n14383 ;
  assign n19377 = x[66] & n12631 ;
  assign n19378 = n19376 | n19377 ;
  assign n19379 = n12700 | n19378 ;
  assign n27910 = ~n19379 ;
  assign n19380 = x[11] & n27910 ;
  assign n19381 = n27892 & n19379 ;
  assign n19382 = n19380 | n19381 ;
  assign n19383 = n19375 & n19382 ;
  assign n19397 = n19375 | n19382 ;
  assign n27911 = ~n19383 ;
  assign n20697 = n27911 & n19397 ;
  assign n15315 = n6379 & n15308 ;
  assign n15287 = x[67] & n15246 ;
  assign n17275 = x[68] & n16288 ;
  assign n20698 = n15287 | n17275 ;
  assign n20699 = x[69] & n15244 ;
  assign n20700 = n20698 | n20699 ;
  assign n20701 = n15315 | n20700 ;
  assign n27912 = ~n20701 ;
  assign n20702 = x[8] & n27912 ;
  assign n20703 = n27845 & n20701 ;
  assign n20704 = n20702 | n20703 ;
  assign n27913 = ~n20704 ;
  assign n20705 = n20697 & n27913 ;
  assign n27914 = ~n20697 ;
  assign n20753 = n27914 & n20704 ;
  assign n20754 = n20705 | n20753 ;
  assign n21161 = n20715 | n21160 ;
  assign n21162 = n20754 | n21161 ;
  assign n21163 = n20754 & n21161 ;
  assign n27915 = ~n21163 ;
  assign n21744 = n21162 & n27915 ;
  assign n27916 = ~n21743 ;
  assign n21845 = n27916 & n21744 ;
  assign n27917 = ~n21744 ;
  assign n21846 = n21743 & n27917 ;
  assign n21847 = n21845 | n21846 ;
  assign n27918 = ~n21752 ;
  assign n21756 = n27918 & n21754 ;
  assign n27919 = ~n21754 ;
  assign n22136 = n21752 & n27919 ;
  assign n22137 = n21756 | n22136 ;
  assign n22160 = n22137 & n22158 ;
  assign n22161 = n21755 | n22160 ;
  assign n27920 = ~n21847 ;
  assign n22162 = n27920 & n22161 ;
  assign n27921 = ~n22161 ;
  assign n22831 = n21847 & n27921 ;
  assign n22832 = n22162 | n22831 ;
  assign n486 = n484 & n485 ;
  assign n487 = n26995 | n486 ;
  assign n27649 = x[74] & x[75] ;
  assign n488 = x[74] | x[75] ;
  assign n27922 = ~n27649 ;
  assign n3286 = n27922 & n488 ;
  assign n3287 = n487 | n3286 ;
  assign n3288 = n487 & n3286 ;
  assign n27923 = ~n3288 ;
  assign n3289 = n3287 & n27923 ;
  assign n19657 = n3289 & n19656 ;
  assign n19779 = x[73] & n19723 ;
  assign n19833 = x[74] & n19829 ;
  assign n22833 = n19779 | n19833 ;
  assign n22834 = x[75] & n19655 ;
  assign n22835 = n22833 | n22834 ;
  assign n22836 = n19657 | n22835 ;
  assign n27924 = ~n22836 ;
  assign n22837 = x[2] & n27924 ;
  assign n22838 = n27790 & n22836 ;
  assign n22839 = n22837 | n22838 ;
  assign n27925 = ~n22839 ;
  assign n22840 = n22832 & n27925 ;
  assign n27926 = ~n22832 ;
  assign n22841 = n27926 & n22839 ;
  assign n22842 = n22840 | n22841 ;
  assign n22843 = n22830 | n22842 ;
  assign n22845 = n22830 & n22842 ;
  assign n27927 = ~n22845 ;
  assign n140 = n22843 & n27927 ;
  assign n489 = n487 & n488 ;
  assign n490 = n27649 | n489 ;
  assign n26915 = x[75] & x[76] ;
  assign n491 = x[75] | x[76] ;
  assign n27928 = ~n26915 ;
  assign n2747 = n27928 & n491 ;
  assign n2748 = n490 & n2747 ;
  assign n2749 = n490 | n2747 ;
  assign n27929 = ~n2748 ;
  assign n2750 = n27929 & n2749 ;
  assign n19680 = n2750 & n19656 ;
  assign n19759 = x[74] & n19723 ;
  assign n19869 = x[75] & n19829 ;
  assign n22688 = n19759 | n19869 ;
  assign n22689 = x[76] & n19655 ;
  assign n22690 = n22688 | n22689 ;
  assign n22691 = n19680 | n22690 ;
  assign n22692 = x[2] | n22691 ;
  assign n22693 = x[2] & n22691 ;
  assign n27930 = ~n22693 ;
  assign n22694 = n22692 & n27930 ;
  assign n15337 = n5976 & n15308 ;
  assign n15254 = x[68] & n15246 ;
  assign n17288 = x[69] & n16288 ;
  assign n20682 = n15254 | n17288 ;
  assign n20683 = x[70] & n15244 ;
  assign n20684 = n20682 | n20683 ;
  assign n20685 = n15337 | n20684 ;
  assign n27931 = ~n20685 ;
  assign n20686 = x[8] & n27931 ;
  assign n20687 = n27845 & n20685 ;
  assign n20688 = n20686 | n20687 ;
  assign n12728 = n6494 & n12695 ;
  assign n12694 = x[65] & n12633 ;
  assign n14409 = x[66] & n13533 ;
  assign n19388 = n12694 | n14409 ;
  assign n19389 = x[67] & n12631 ;
  assign n19390 = n19388 | n19389 ;
  assign n19391 = n12728 | n19390 ;
  assign n27932 = ~n19391 ;
  assign n19392 = x[11] & n27932 ;
  assign n19393 = n27892 & n19391 ;
  assign n19394 = n19392 | n19393 ;
  assign n267 = x[11] & x[12] ;
  assign n10475 = x[11] | x[12] ;
  assign n27933 = ~n267 ;
  assign n10476 = n27933 & n10475 ;
  assign n18088 = x[64] & n10476 ;
  assign n27934 = ~n18088 ;
  assign n19385 = n27934 & n19383 ;
  assign n20340 = n18088 & n27911 ;
  assign n20341 = n19385 | n20340 ;
  assign n20342 = n19394 | n20341 ;
  assign n20343 = n19394 & n20341 ;
  assign n27935 = ~n20343 ;
  assign n20692 = n20342 & n27935 ;
  assign n27936 = ~n20688 ;
  assign n20693 = n27936 & n20692 ;
  assign n27937 = ~n20692 ;
  assign n20695 = n20688 & n27937 ;
  assign n20696 = n20693 | n20695 ;
  assign n20706 = n20697 & n20704 ;
  assign n20746 = n20738 & n20745 ;
  assign n20749 = n20735 | n20746 ;
  assign n20751 = n20749 & n20750 ;
  assign n20752 = n20715 | n20751 ;
  assign n20755 = n20752 & n20754 ;
  assign n20756 = n20706 | n20755 ;
  assign n20757 = n20696 | n20756 ;
  assign n20758 = n20696 & n20756 ;
  assign n27938 = ~n20758 ;
  assign n21724 = n20757 & n27938 ;
  assign n18442 = n3733 & n18392 ;
  assign n18372 = x[71] & n18329 ;
  assign n18519 = x[72] & n18514 ;
  assign n21725 = n18372 | n18519 ;
  assign n21726 = x[73] & n18327 ;
  assign n21727 = n21725 | n21726 ;
  assign n21728 = n18442 | n21727 ;
  assign n27939 = ~n21728 ;
  assign n21729 = x[5] & n27939 ;
  assign n21730 = n27813 & n21728 ;
  assign n21731 = n21729 | n21730 ;
  assign n27940 = ~n21731 ;
  assign n21732 = n21724 & n27940 ;
  assign n27941 = ~n21724 ;
  assign n22134 = n27941 & n21731 ;
  assign n22135 = n21732 | n22134 ;
  assign n21745 = n21743 & n21744 ;
  assign n22163 = n21743 | n21744 ;
  assign n27942 = ~n21745 ;
  assign n22164 = n27942 & n22163 ;
  assign n22165 = n22161 & n22164 ;
  assign n22166 = n21745 | n22165 ;
  assign n22167 = n22135 | n22166 ;
  assign n22168 = n22135 & n22166 ;
  assign n27943 = ~n22168 ;
  assign n22695 = n22167 & n27943 ;
  assign n22696 = n22694 & n22695 ;
  assign n22697 = n22694 | n22695 ;
  assign n27944 = ~n22696 ;
  assign n22698 = n27944 & n22697 ;
  assign n22844 = n22832 & n22839 ;
  assign n22846 = n22844 | n22845 ;
  assign n22847 = n22698 & n22846 ;
  assign n27635 = n22698 | n22846 ;
  assign n27945 = ~n22847 ;
  assign n141 = n27945 & n27635 ;
  assign n22848 = n22696 | n22847 ;
  assign n20694 = n20688 & n20692 ;
  assign n21151 = n20688 | n20692 ;
  assign n27946 = ~n20694 ;
  assign n21152 = n27946 & n21151 ;
  assign n27947 = ~n20756 ;
  assign n21153 = n27947 & n21152 ;
  assign n27948 = ~n21152 ;
  assign n21734 = n20756 & n27948 ;
  assign n21735 = n21153 | n21734 ;
  assign n22133 = n21731 & n21735 ;
  assign n22169 = n22133 | n22168 ;
  assign n15309 = n4790 & n15308 ;
  assign n15247 = x[69] & n15246 ;
  assign n17277 = x[70] & n16288 ;
  assign n20669 = n15247 | n17277 ;
  assign n20670 = x[71] & n15244 ;
  assign n20671 = n20669 | n20670 ;
  assign n20672 = n15309 | n20671 ;
  assign n27949 = ~n20672 ;
  assign n20673 = x[8] & n27949 ;
  assign n20674 = n27845 & n20672 ;
  assign n20675 = n20673 | n20674 ;
  assign n19384 = n18088 & n19383 ;
  assign n20344 = n19384 | n20343 ;
  assign n12758 = n6408 & n12695 ;
  assign n12645 = x[66] & n12633 ;
  assign n14350 = x[67] & n13533 ;
  assign n19356 = n12645 | n14350 ;
  assign n19357 = x[68] & n12631 ;
  assign n19358 = n19356 | n19357 ;
  assign n19359 = n12758 | n19358 ;
  assign n27950 = ~n19359 ;
  assign n19360 = x[11] & n27950 ;
  assign n19361 = n27892 & n19359 ;
  assign n19362 = n19360 | n19361 ;
  assign n18089 = x[14] & n27934 ;
  assign n268 = x[13] & x[14] ;
  assign n10477 = x[13] | x[14] ;
  assign n27951 = ~n268 ;
  assign n10478 = n27951 & n10477 ;
  assign n10542 = n10476 & n10478 ;
  assign n10585 = n6437 & n10542 ;
  assign n266 = x[12] & x[13] ;
  assign n10473 = x[12] | x[13] ;
  assign n27952 = ~n266 ;
  assign n10474 = n27952 & n10473 ;
  assign n27953 = ~n10476 ;
  assign n11232 = n10474 & n27953 ;
  assign n18090 = x[64] & n11232 ;
  assign n27954 = ~n10478 ;
  assign n10479 = n10476 & n27954 ;
  assign n18091 = x[65] & n10479 ;
  assign n18092 = n18090 | n18091 ;
  assign n18093 = n10585 | n18092 ;
  assign n27955 = ~n18093 ;
  assign n18094 = x[14] & n27955 ;
  assign n27956 = ~x[14] ;
  assign n18095 = n27956 & n18093 ;
  assign n18096 = n18094 | n18095 ;
  assign n18097 = n18089 | n18096 ;
  assign n18098 = n18089 & n18096 ;
  assign n27957 = ~n18098 ;
  assign n19363 = n18097 & n27957 ;
  assign n19364 = n19362 & n19363 ;
  assign n19399 = n19362 | n19363 ;
  assign n27958 = ~n19364 ;
  assign n20345 = n27958 & n19399 ;
  assign n20346 = n20344 & n20345 ;
  assign n20676 = n20344 | n20345 ;
  assign n27959 = ~n20346 ;
  assign n20677 = n27959 & n20676 ;
  assign n20678 = n20675 & n20677 ;
  assign n20680 = n20675 | n20677 ;
  assign n27960 = ~n20678 ;
  assign n20681 = n27960 & n20680 ;
  assign n19386 = n18088 | n19383 ;
  assign n27961 = ~n19384 ;
  assign n19387 = n27961 & n19386 ;
  assign n27962 = ~n19394 ;
  assign n19396 = n19387 & n27962 ;
  assign n27963 = ~n19387 ;
  assign n20689 = n27963 & n19394 ;
  assign n20690 = n19396 | n20689 ;
  assign n20691 = n20688 & n20690 ;
  assign n21164 = n20706 | n21163 ;
  assign n21165 = n21152 & n21164 ;
  assign n21166 = n20691 | n21165 ;
  assign n27964 = ~n21166 ;
  assign n21167 = n20681 & n27964 ;
  assign n27965 = ~n20681 ;
  assign n21714 = n27965 & n21166 ;
  assign n21715 = n21167 | n21714 ;
  assign n18395 = n2722 & n18392 ;
  assign n18362 = x[72] & n18329 ;
  assign n18556 = x[73] & n18514 ;
  assign n21716 = n18362 | n18556 ;
  assign n21717 = x[74] & n18327 ;
  assign n21718 = n21716 | n21717 ;
  assign n21719 = n18395 | n21718 ;
  assign n27966 = ~n21719 ;
  assign n21720 = x[5] & n27966 ;
  assign n21721 = n27813 & n21719 ;
  assign n21722 = n21720 | n21721 ;
  assign n21852 = n21715 | n21722 ;
  assign n27967 = ~n20675 ;
  assign n20679 = n27967 & n20677 ;
  assign n27968 = ~n20677 ;
  assign n21149 = n20675 & n27968 ;
  assign n21150 = n20679 | n21149 ;
  assign n21168 = n21150 | n21166 ;
  assign n21169 = n21150 & n21166 ;
  assign n27969 = ~n21169 ;
  assign n22131 = n21168 & n27969 ;
  assign n22132 = n21722 & n22131 ;
  assign n27970 = ~n22132 ;
  assign n22849 = n21852 & n27970 ;
  assign n27971 = ~n22849 ;
  assign n22850 = n22169 & n27971 ;
  assign n21723 = n21715 & n21722 ;
  assign n21733 = n21724 & n21731 ;
  assign n21736 = n21731 | n21735 ;
  assign n21842 = n21768 | n21841 ;
  assign n21843 = n21758 & n21842 ;
  assign n21844 = n21755 | n21843 ;
  assign n21848 = n21844 & n21847 ;
  assign n21849 = n21745 | n21848 ;
  assign n21850 = n21736 & n21849 ;
  assign n21851 = n21733 | n21850 ;
  assign n21853 = n21851 & n21852 ;
  assign n21854 = n21723 | n21853 ;
  assign n27972 = ~n21854 ;
  assign n22851 = n21852 & n27972 ;
  assign n22852 = n22850 | n22851 ;
  assign n492 = n490 & n491 ;
  assign n493 = n26915 | n492 ;
  assign n27647 = x[76] & x[77] ;
  assign n494 = x[76] | x[77] ;
  assign n27973 = ~n27647 ;
  assign n1772 = n27973 & n494 ;
  assign n1773 = n493 | n1772 ;
  assign n1774 = n493 & n1772 ;
  assign n27974 = ~n1774 ;
  assign n1775 = n1773 & n27974 ;
  assign n19689 = n1775 & n19656 ;
  assign n19729 = x[75] & n19723 ;
  assign n19856 = x[76] & n19829 ;
  assign n22853 = n19729 | n19856 ;
  assign n22854 = x[77] & n19655 ;
  assign n22855 = n22853 | n22854 ;
  assign n22856 = n19689 | n22855 ;
  assign n27975 = ~n22856 ;
  assign n22857 = x[2] & n27975 ;
  assign n22858 = n27790 & n22856 ;
  assign n22859 = n22857 | n22858 ;
  assign n27976 = ~n22859 ;
  assign n22860 = n22852 & n27976 ;
  assign n27977 = ~n22852 ;
  assign n22861 = n27977 & n22859 ;
  assign n22862 = n22860 | n22861 ;
  assign n22863 = n22848 | n22862 ;
  assign n22865 = n22848 & n22862 ;
  assign n27978 = ~n22865 ;
  assign n142 = n22863 & n27978 ;
  assign n22864 = n22852 & n22859 ;
  assign n22866 = n22864 | n22865 ;
  assign n495 = n493 & n494 ;
  assign n496 = n27647 | n495 ;
  assign n26823 = x[77] & x[78] ;
  assign n497 = x[77] | x[78] ;
  assign n27979 = ~n26823 ;
  assign n2081 = n27979 & n497 ;
  assign n2082 = n496 & n2081 ;
  assign n2083 = n496 | n2081 ;
  assign n27980 = ~n2082 ;
  assign n2084 = n27980 & n2083 ;
  assign n19701 = n2084 & n19656 ;
  assign n19732 = x[76] & n19723 ;
  assign n19877 = x[77] & n19829 ;
  assign n22867 = n19732 | n19877 ;
  assign n22868 = x[78] & n19655 ;
  assign n22869 = n22867 | n22868 ;
  assign n22870 = n19701 | n22869 ;
  assign n22871 = x[2] | n22870 ;
  assign n22872 = x[2] & n22870 ;
  assign n27981 = ~n22872 ;
  assign n22873 = n22871 & n27981 ;
  assign n18398 = n3289 & n18392 ;
  assign n18373 = x[73] & n18329 ;
  assign n18521 = x[74] & n18514 ;
  assign n21704 = n18373 | n18521 ;
  assign n21705 = x[75] & n18327 ;
  assign n21706 = n21704 | n21705 ;
  assign n21707 = n18398 | n21706 ;
  assign n27982 = ~n21707 ;
  assign n21708 = x[5] & n27982 ;
  assign n21709 = n27813 & n21707 ;
  assign n21710 = n21708 | n21709 ;
  assign n21170 = n20678 | n21169 ;
  assign n10544 = n6466 & n10542 ;
  assign n10480 = n27953 & n10478 ;
  assign n27983 = ~n10474 ;
  assign n10481 = n27983 & n10480 ;
  assign n10505 = x[64] & n10481 ;
  assign n11885 = x[65] & n11232 ;
  assign n18099 = n10505 | n11885 ;
  assign n18100 = x[66] & n10479 ;
  assign n18101 = n18099 | n18100 ;
  assign n18102 = n10544 | n18101 ;
  assign n27984 = ~n18102 ;
  assign n18103 = x[14] & n27984 ;
  assign n18104 = n27956 & n18102 ;
  assign n18105 = n18103 | n18104 ;
  assign n18106 = n18098 & n18105 ;
  assign n18120 = n18098 | n18105 ;
  assign n27985 = ~n18106 ;
  assign n19347 = n27985 & n18120 ;
  assign n12757 = n6379 & n12695 ;
  assign n12638 = x[67] & n12633 ;
  assign n14387 = x[68] & n13533 ;
  assign n19348 = n12638 | n14387 ;
  assign n19349 = x[69] & n12631 ;
  assign n19350 = n19348 | n19349 ;
  assign n19351 = n12757 | n19350 ;
  assign n27986 = ~n19351 ;
  assign n19352 = x[11] & n27986 ;
  assign n19353 = n27892 & n19351 ;
  assign n19354 = n19352 | n19353 ;
  assign n19402 = n19347 | n19354 ;
  assign n19355 = n19347 & n19354 ;
  assign n19395 = n19387 & n19394 ;
  assign n19398 = n19384 | n19395 ;
  assign n19400 = n19398 & n19399 ;
  assign n19401 = n19364 | n19400 ;
  assign n19403 = n19401 & n19402 ;
  assign n19405 = n19355 | n19403 ;
  assign n27987 = ~n19405 ;
  assign n19406 = n19402 & n27987 ;
  assign n27988 = ~n19355 ;
  assign n19404 = n27988 & n19402 ;
  assign n20347 = n19364 | n20346 ;
  assign n27989 = ~n19404 ;
  assign n20658 = n27989 & n20347 ;
  assign n20659 = n19406 | n20658 ;
  assign n15317 = n3701 & n15308 ;
  assign n15248 = x[70] & n15246 ;
  assign n17278 = x[71] & n16288 ;
  assign n20660 = n15248 | n17278 ;
  assign n20661 = x[72] & n15244 ;
  assign n20662 = n20660 | n20661 ;
  assign n20663 = n15317 | n20662 ;
  assign n27990 = ~n20663 ;
  assign n20664 = x[8] & n27990 ;
  assign n20665 = n27845 & n20663 ;
  assign n20666 = n20664 | n20665 ;
  assign n20667 = n20659 | n20666 ;
  assign n20668 = n20659 & n20666 ;
  assign n27991 = ~n20668 ;
  assign n21171 = n20667 & n27991 ;
  assign n21172 = n21170 & n21171 ;
  assign n21711 = n21170 | n21171 ;
  assign n27992 = ~n21172 ;
  assign n21712 = n27992 & n21711 ;
  assign n21713 = n21710 & n21712 ;
  assign n21855 = n21710 | n21712 ;
  assign n27993 = ~n21713 ;
  assign n21856 = n27993 & n21855 ;
  assign n22170 = n21722 | n22131 ;
  assign n22171 = n22169 & n22170 ;
  assign n22172 = n22132 | n22171 ;
  assign n27994 = ~n22172 ;
  assign n22173 = n21856 & n27994 ;
  assign n27995 = ~n21856 ;
  assign n22874 = n27995 & n22172 ;
  assign n22875 = n22173 | n22874 ;
  assign n27996 = ~n22875 ;
  assign n22876 = n22873 & n27996 ;
  assign n27997 = ~n22873 ;
  assign n22877 = n27997 & n22875 ;
  assign n22878 = n22876 | n22877 ;
  assign n22879 = n22866 & n22878 ;
  assign n27638 = n22866 | n22878 ;
  assign n27998 = ~n22879 ;
  assign n143 = n27998 & n27638 ;
  assign n22880 = n22873 & n22875 ;
  assign n22881 = n22879 | n22880 ;
  assign n498 = n496 & n497 ;
  assign n499 = n26823 | n498 ;
  assign n27646 = x[78] & x[79] ;
  assign n500 = x[78] | x[79] ;
  assign n27999 = ~n27646 ;
  assign n1738 = n27999 & n500 ;
  assign n1739 = n499 | n1738 ;
  assign n1740 = n499 & n1738 ;
  assign n28000 = ~n1740 ;
  assign n1741 = n1739 & n28000 ;
  assign n19663 = n1741 & n19656 ;
  assign n19730 = x[77] & n19723 ;
  assign n19840 = x[78] & n19829 ;
  assign n22675 = n19730 | n19840 ;
  assign n22676 = x[79] & n19655 ;
  assign n22677 = n22675 | n22676 ;
  assign n22678 = n19663 | n22677 ;
  assign n28001 = ~n22678 ;
  assign n22679 = x[2] & n28001 ;
  assign n22680 = n27790 & n22678 ;
  assign n22681 = n22679 | n22680 ;
  assign n21857 = n21854 & n21856 ;
  assign n21858 = n21713 | n21857 ;
  assign n18406 = n2750 & n18392 ;
  assign n18367 = x[74] & n18329 ;
  assign n18557 = x[75] & n18514 ;
  assign n21691 = n18367 | n18557 ;
  assign n21692 = x[76] & n18327 ;
  assign n21693 = n21691 | n21692 ;
  assign n21694 = n18406 | n21693 ;
  assign n28002 = ~n21694 ;
  assign n21695 = x[5] & n28002 ;
  assign n21696 = n27813 & n21694 ;
  assign n21697 = n21695 | n21696 ;
  assign n12696 = n5976 & n12695 ;
  assign n12634 = x[68] & n12633 ;
  assign n14392 = x[69] & n13533 ;
  assign n19337 = n12634 | n14392 ;
  assign n19338 = x[70] & n12631 ;
  assign n19339 = n19337 | n19338 ;
  assign n19340 = n12696 | n19339 ;
  assign n28003 = ~n19340 ;
  assign n19341 = x[11] & n28003 ;
  assign n19342 = n27892 & n19340 ;
  assign n19343 = n19341 | n19342 ;
  assign n10604 = n6494 & n10542 ;
  assign n10541 = x[65] & n10481 ;
  assign n11919 = x[66] & n11232 ;
  assign n18111 = n10541 | n11919 ;
  assign n18112 = x[67] & n10479 ;
  assign n18113 = n18111 | n18112 ;
  assign n18114 = n10604 | n18113 ;
  assign n28004 = ~n18114 ;
  assign n18115 = x[14] & n28004 ;
  assign n18116 = n27956 & n18114 ;
  assign n18117 = n18115 | n18116 ;
  assign n264 = x[14] & x[15] ;
  assign n8639 = x[14] | x[15] ;
  assign n28005 = ~n264 ;
  assign n8640 = n28005 & n8639 ;
  assign n17014 = x[64] & n8640 ;
  assign n28006 = ~n17014 ;
  assign n18108 = n28006 & n18106 ;
  assign n19073 = n17014 & n27985 ;
  assign n19074 = n18108 | n19073 ;
  assign n19075 = n18117 | n19074 ;
  assign n19076 = n18117 & n19074 ;
  assign n28007 = ~n19076 ;
  assign n19407 = n19075 & n28007 ;
  assign n28008 = ~n19343 ;
  assign n19408 = n28008 & n19407 ;
  assign n28009 = ~n19407 ;
  assign n19410 = n19343 & n28009 ;
  assign n19411 = n19408 | n19410 ;
  assign n20348 = n19402 & n20347 ;
  assign n20349 = n19355 | n20348 ;
  assign n28010 = ~n19411 ;
  assign n20350 = n28010 & n20349 ;
  assign n28011 = ~n20349 ;
  assign n20655 = n19411 & n28011 ;
  assign n20656 = n20350 | n20655 ;
  assign n15310 = n3733 & n15308 ;
  assign n15266 = x[71] & n15246 ;
  assign n17299 = x[72] & n16288 ;
  assign n20647 = n15266 | n17299 ;
  assign n20648 = x[73] & n15244 ;
  assign n20649 = n20647 | n20648 ;
  assign n20650 = n15310 | n20649 ;
  assign n28012 = ~n20650 ;
  assign n20652 = x[8] & n28012 ;
  assign n20764 = n27845 & n20650 ;
  assign n20765 = n20652 | n20764 ;
  assign n28013 = ~n20656 ;
  assign n20766 = n28013 & n20765 ;
  assign n28014 = ~n20765 ;
  assign n20767 = n20656 & n28014 ;
  assign n20768 = n20766 | n20767 ;
  assign n21173 = n20668 | n21172 ;
  assign n21174 = n20768 & n21173 ;
  assign n21698 = n20767 | n21173 ;
  assign n21699 = n20766 | n21698 ;
  assign n28015 = ~n21174 ;
  assign n21700 = n28015 & n21699 ;
  assign n28016 = ~n21700 ;
  assign n21701 = n21697 & n28016 ;
  assign n28017 = ~n21697 ;
  assign n21859 = n28017 & n21700 ;
  assign n21860 = n21701 | n21859 ;
  assign n21861 = n21858 & n21860 ;
  assign n21703 = n21697 & n21700 ;
  assign n28018 = ~n21703 ;
  assign n22682 = n21700 & n28018 ;
  assign n22683 = n21858 | n22682 ;
  assign n22684 = n21701 | n22683 ;
  assign n28019 = ~n21861 ;
  assign n22685 = n28019 & n22684 ;
  assign n22686 = n22681 | n22685 ;
  assign n22687 = n22681 & n22685 ;
  assign n28020 = ~n22687 ;
  assign n22882 = n22686 & n28020 ;
  assign n22883 = n22881 & n22882 ;
  assign n28021 = ~n22685 ;
  assign n27640 = n22681 & n28021 ;
  assign n28022 = ~n22681 ;
  assign n27641 = n28022 & n22685 ;
  assign n27642 = n22881 | n27641 ;
  assign n27643 = n27640 | n27642 ;
  assign n28023 = ~n22883 ;
  assign n144 = n28023 & n27643 ;
  assign n22884 = n22687 | n22883 ;
  assign n501 = n499 & n500 ;
  assign n502 = n27646 | n501 ;
  assign n26737 = x[79] & x[80] ;
  assign n503 = x[79] | x[80] ;
  assign n28024 = ~n26737 ;
  assign n1267 = n28024 & n503 ;
  assign n1268 = n502 & n1267 ;
  assign n1269 = n502 | n1267 ;
  assign n28025 = ~n1268 ;
  assign n1270 = n28025 & n1269 ;
  assign n19674 = n1270 & n19656 ;
  assign n19761 = x[78] & n19723 ;
  assign n19832 = x[79] & n19829 ;
  assign n22885 = n19761 | n19832 ;
  assign n22886 = x[80] & n19655 ;
  assign n22887 = n22885 | n22886 ;
  assign n22888 = n19674 | n22887 ;
  assign n22889 = x[2] | n22888 ;
  assign n22890 = x[2] & n22888 ;
  assign n28026 = ~n22890 ;
  assign n22891 = n22889 & n28026 ;
  assign n21862 = n21703 | n21861 ;
  assign n18401 = n1775 & n18392 ;
  assign n18335 = x[75] & n18329 ;
  assign n18522 = x[76] & n18514 ;
  assign n21681 = n18335 | n18522 ;
  assign n21682 = x[77] & n18327 ;
  assign n21683 = n21681 | n21682 ;
  assign n21684 = n18401 | n21683 ;
  assign n28027 = ~n21684 ;
  assign n21685 = x[5] & n28027 ;
  assign n21686 = n27813 & n21684 ;
  assign n21687 = n21685 | n21686 ;
  assign n21148 = n20656 & n20765 ;
  assign n21175 = n21148 | n21174 ;
  assign n15312 = n2722 & n15308 ;
  assign n15249 = x[72] & n15246 ;
  assign n17281 = x[73] & n16288 ;
  assign n20637 = n15249 | n17281 ;
  assign n20638 = x[74] & n15244 ;
  assign n20639 = n20637 | n20638 ;
  assign n20640 = n15312 | n20639 ;
  assign n28028 = ~n20640 ;
  assign n20641 = x[8] & n28028 ;
  assign n20642 = n27845 & n20640 ;
  assign n20643 = n20641 | n20642 ;
  assign n18107 = n17014 & n18106 ;
  assign n18109 = n17014 | n18106 ;
  assign n28029 = ~n18107 ;
  assign n18110 = n28029 & n18109 ;
  assign n28030 = ~n18117 ;
  assign n18119 = n18110 & n28030 ;
  assign n28031 = ~n18110 ;
  assign n19344 = n28031 & n18117 ;
  assign n19345 = n18119 | n19344 ;
  assign n19346 = n19343 & n19345 ;
  assign n19412 = n19405 & n19411 ;
  assign n19413 = n19346 | n19412 ;
  assign n12704 = n4790 & n12695 ;
  assign n12635 = x[69] & n12633 ;
  assign n14353 = x[70] & n13533 ;
  assign n19327 = n12635 | n14353 ;
  assign n19328 = x[71] & n12631 ;
  assign n19329 = n19327 | n19328 ;
  assign n19330 = n12704 | n19329 ;
  assign n28032 = ~n19330 ;
  assign n19331 = x[11] & n28032 ;
  assign n19332 = n27892 & n19330 ;
  assign n19333 = n19331 | n19332 ;
  assign n19077 = n18107 | n19076 ;
  assign n10603 = n6408 & n10542 ;
  assign n10501 = x[66] & n10481 ;
  assign n11927 = x[67] & n11232 ;
  assign n18079 = n10501 | n11927 ;
  assign n18080 = x[68] & n10479 ;
  assign n18081 = n18079 | n18080 ;
  assign n18082 = n10603 | n18081 ;
  assign n28033 = ~n18082 ;
  assign n18083 = x[14] & n28033 ;
  assign n18084 = n27956 & n18082 ;
  assign n18085 = n18083 | n18084 ;
  assign n17015 = x[17] & n28006 ;
  assign n265 = x[16] & x[17] ;
  assign n8641 = x[16] | x[17] ;
  assign n28034 = ~n265 ;
  assign n8642 = n28034 & n8641 ;
  assign n8706 = n8640 & n8642 ;
  assign n8757 = n6437 & n8706 ;
  assign n263 = x[15] & x[16] ;
  assign n8637 = x[15] | x[16] ;
  assign n28035 = ~n263 ;
  assign n8638 = n28035 & n8637 ;
  assign n28036 = ~n8640 ;
  assign n9278 = n8638 & n28036 ;
  assign n17016 = x[64] & n9278 ;
  assign n28037 = ~n8642 ;
  assign n8643 = n8640 & n28037 ;
  assign n17017 = x[65] & n8643 ;
  assign n17018 = n17016 | n17017 ;
  assign n17019 = n8757 | n17018 ;
  assign n28038 = ~n17019 ;
  assign n17020 = x[17] & n28038 ;
  assign n28039 = ~x[17] ;
  assign n17021 = n28039 & n17019 ;
  assign n17022 = n17020 | n17021 ;
  assign n17023 = n17015 | n17022 ;
  assign n17024 = n17015 & n17022 ;
  assign n28040 = ~n17024 ;
  assign n18086 = n17023 & n28040 ;
  assign n18087 = n18085 & n18086 ;
  assign n18122 = n18085 | n18086 ;
  assign n28041 = ~n18087 ;
  assign n19078 = n28041 & n18122 ;
  assign n19079 = n19077 & n19078 ;
  assign n19334 = n19077 | n19078 ;
  assign n28042 = ~n19079 ;
  assign n19335 = n28042 & n19334 ;
  assign n19336 = n19333 & n19335 ;
  assign n19414 = n19333 | n19335 ;
  assign n28043 = ~n19336 ;
  assign n19415 = n28043 & n19414 ;
  assign n19416 = n19413 & n19415 ;
  assign n20644 = n19413 | n19415 ;
  assign n28044 = ~n19416 ;
  assign n20645 = n28044 & n20644 ;
  assign n20646 = n20643 & n20645 ;
  assign n20771 = n20643 | n20645 ;
  assign n28045 = ~n20646 ;
  assign n21176 = n28045 & n20771 ;
  assign n21177 = n21175 & n21176 ;
  assign n21688 = n21175 | n21176 ;
  assign n28046 = ~n21177 ;
  assign n21689 = n28046 & n21688 ;
  assign n21690 = n21687 & n21689 ;
  assign n21863 = n21687 | n21689 ;
  assign n28047 = ~n21690 ;
  assign n21864 = n28047 & n21863 ;
  assign n21865 = n21862 & n21864 ;
  assign n22892 = n21862 | n21864 ;
  assign n28048 = ~n21865 ;
  assign n22893 = n28048 & n22892 ;
  assign n22894 = n22891 & n22893 ;
  assign n22895 = n22891 | n22893 ;
  assign n28049 = ~n22894 ;
  assign n22896 = n28049 & n22895 ;
  assign n22897 = n22884 & n22896 ;
  assign n27645 = n22884 | n22896 ;
  assign n28050 = ~n22897 ;
  assign n145 = n28050 & n27645 ;
  assign n504 = n502 & n503 ;
  assign n505 = n26737 | n504 ;
  assign n27644 = x[80] & x[81] ;
  assign n506 = x[80] | x[81] ;
  assign n28051 = ~n27644 ;
  assign n1026 = n28051 & n506 ;
  assign n28052 = ~n505 ;
  assign n1027 = n28052 & n1026 ;
  assign n28053 = ~n1026 ;
  assign n1028 = n505 & n28053 ;
  assign n1029 = n1027 | n1028 ;
  assign n19668 = n1029 & n19656 ;
  assign n19767 = x[79] & n19723 ;
  assign n19837 = x[80] & n19829 ;
  assign n22663 = n19767 | n19837 ;
  assign n22664 = x[81] & n19655 ;
  assign n22665 = n22663 | n22664 ;
  assign n22666 = n19668 | n22665 ;
  assign n28054 = ~n22666 ;
  assign n22667 = x[2] & n28054 ;
  assign n22668 = n27790 & n22666 ;
  assign n22669 = n22667 | n22668 ;
  assign n21866 = n21690 | n21865 ;
  assign n18402 = n2084 & n18392 ;
  assign n18331 = x[76] & n18329 ;
  assign n18536 = x[77] & n18514 ;
  assign n21671 = n18331 | n18536 ;
  assign n21672 = x[78] & n18327 ;
  assign n21673 = n21671 | n21672 ;
  assign n21674 = n18402 | n21673 ;
  assign n28055 = ~n21674 ;
  assign n21675 = x[5] & n28055 ;
  assign n21676 = n27813 & n21674 ;
  assign n21677 = n21675 | n21676 ;
  assign n15336 = n3289 & n15308 ;
  assign n15269 = x[73] & n15246 ;
  assign n17331 = x[74] & n16288 ;
  assign n20627 = n15269 | n17331 ;
  assign n20628 = x[75] & n15244 ;
  assign n20629 = n20627 | n20628 ;
  assign n20630 = n15336 | n20629 ;
  assign n28056 = ~n20630 ;
  assign n20631 = x[8] & n28056 ;
  assign n20632 = n27845 & n20630 ;
  assign n20633 = n20631 | n20632 ;
  assign n19417 = n19336 | n19416 ;
  assign n8715 = n6466 & n8706 ;
  assign n8644 = n28036 & n8642 ;
  assign n28057 = ~n8638 ;
  assign n8645 = n28057 & n8644 ;
  assign n8646 = x[64] & n8645 ;
  assign n9865 = x[65] & n9278 ;
  assign n17025 = n8646 | n9865 ;
  assign n17026 = x[66] & n8643 ;
  assign n17027 = n17025 | n17026 ;
  assign n17028 = n8715 | n17027 ;
  assign n28058 = ~n17028 ;
  assign n17029 = x[17] & n28058 ;
  assign n17030 = n28039 & n17028 ;
  assign n17031 = n17029 | n17030 ;
  assign n17032 = n17024 | n17031 ;
  assign n17033 = n17024 & n17031 ;
  assign n28059 = ~n17033 ;
  assign n18070 = n17032 & n28059 ;
  assign n10593 = n6379 & n10542 ;
  assign n10482 = x[67] & n10481 ;
  assign n11928 = x[68] & n11232 ;
  assign n18071 = n10482 | n11928 ;
  assign n18072 = x[69] & n10479 ;
  assign n18073 = n18071 | n18072 ;
  assign n18074 = n10593 | n18073 ;
  assign n28060 = ~n18074 ;
  assign n18075 = x[14] & n28060 ;
  assign n18076 = n27956 & n18074 ;
  assign n18077 = n18075 | n18076 ;
  assign n18125 = n18070 | n18077 ;
  assign n18078 = n18070 & n18077 ;
  assign n18118 = n18110 & n18117 ;
  assign n18121 = n18107 | n18118 ;
  assign n18123 = n18121 & n18122 ;
  assign n18124 = n18087 | n18123 ;
  assign n18126 = n18124 & n18125 ;
  assign n18128 = n18078 | n18126 ;
  assign n28061 = ~n18128 ;
  assign n18129 = n18125 & n28061 ;
  assign n28062 = ~n18078 ;
  assign n18127 = n28062 & n18125 ;
  assign n19080 = n18087 | n19079 ;
  assign n28063 = ~n18127 ;
  assign n19316 = n28063 & n19080 ;
  assign n19317 = n18129 | n19316 ;
  assign n12697 = n3701 & n12695 ;
  assign n12646 = x[70] & n12633 ;
  assign n14355 = x[71] & n13533 ;
  assign n19318 = n12646 | n14355 ;
  assign n19319 = x[72] & n12631 ;
  assign n19320 = n19318 | n19319 ;
  assign n19321 = n12697 | n19320 ;
  assign n28064 = ~n19321 ;
  assign n19322 = x[11] & n28064 ;
  assign n19323 = n27892 & n19321 ;
  assign n19324 = n19322 | n19323 ;
  assign n19325 = n19317 | n19324 ;
  assign n19326 = n19317 & n19324 ;
  assign n28065 = ~n19326 ;
  assign n20357 = n19325 & n28065 ;
  assign n28066 = ~n19417 ;
  assign n20359 = n28066 & n20357 ;
  assign n28067 = ~n20357 ;
  assign n20634 = n19417 & n28067 ;
  assign n20635 = n20359 | n20634 ;
  assign n20636 = n20633 & n20635 ;
  assign n20774 = n20633 | n20635 ;
  assign n28068 = ~n20636 ;
  assign n20775 = n28068 & n20774 ;
  assign n21178 = n20646 | n21177 ;
  assign n28069 = ~n21178 ;
  assign n21179 = n20775 & n28069 ;
  assign n28070 = ~n20775 ;
  assign n21678 = n28070 & n21178 ;
  assign n21679 = n21179 | n21678 ;
  assign n21680 = n21677 & n21679 ;
  assign n21867 = n21677 | n21679 ;
  assign n28071 = ~n21680 ;
  assign n22181 = n28071 & n21867 ;
  assign n28072 = ~n21866 ;
  assign n22183 = n28072 & n22181 ;
  assign n28073 = ~n22181 ;
  assign n22670 = n21866 & n28073 ;
  assign n22671 = n22183 | n22670 ;
  assign n22672 = n22669 | n22671 ;
  assign n22673 = n22669 & n22671 ;
  assign n28074 = ~n22673 ;
  assign n22674 = n22672 & n28074 ;
  assign n22898 = n22894 | n22897 ;
  assign n22899 = n22674 | n22898 ;
  assign n22900 = n22674 & n22898 ;
  assign n28075 = ~n22900 ;
  assign n146 = n22899 & n28075 ;
  assign n18410 = n1741 & n18392 ;
  assign n18349 = x[77] & n18329 ;
  assign n18570 = x[78] & n18514 ;
  assign n21661 = n18349 | n18570 ;
  assign n21662 = x[79] & n18327 ;
  assign n21663 = n21661 | n21662 ;
  assign n21664 = n18410 | n21663 ;
  assign n28076 = ~n21664 ;
  assign n21665 = x[5] & n28076 ;
  assign n21666 = n27813 & n21664 ;
  assign n21667 = n21665 | n21666 ;
  assign n20651 = x[8] | n20650 ;
  assign n20653 = x[8] & n20650 ;
  assign n28077 = ~n20653 ;
  assign n20654 = n20651 & n28077 ;
  assign n20657 = n20654 & n20656 ;
  assign n20759 = n20691 | n20758 ;
  assign n20760 = n20681 & n20759 ;
  assign n20761 = n20678 | n20760 ;
  assign n20762 = n20667 & n20761 ;
  assign n20763 = n20668 | n20762 ;
  assign n20769 = n20763 & n20768 ;
  assign n20770 = n20657 | n20769 ;
  assign n20772 = n20770 & n20771 ;
  assign n20773 = n20646 | n20772 ;
  assign n20776 = n20773 & n20775 ;
  assign n20777 = n20636 | n20776 ;
  assign n15332 = n2750 & n15308 ;
  assign n15301 = x[74] & n15246 ;
  assign n17285 = x[75] & n16288 ;
  assign n20617 = n15301 | n17285 ;
  assign n20618 = x[76] & n15244 ;
  assign n20619 = n20617 | n20618 ;
  assign n20620 = n15332 | n20619 ;
  assign n28078 = ~n20620 ;
  assign n20621 = x[8] & n28078 ;
  assign n20622 = n27845 & n20620 ;
  assign n20623 = n20621 | n20622 ;
  assign n10557 = n5976 & n10542 ;
  assign n10483 = x[68] & n10481 ;
  assign n11893 = x[69] & n11232 ;
  assign n18061 = n10483 | n11893 ;
  assign n18062 = x[70] & n10479 ;
  assign n18063 = n18061 | n18062 ;
  assign n18064 = n10557 | n18063 ;
  assign n28079 = ~n18064 ;
  assign n18065 = x[14] & n28079 ;
  assign n18066 = n27956 & n18064 ;
  assign n18067 = n18065 | n18066 ;
  assign n261 = x[17] & x[18] ;
  assign n7094 = x[17] | x[18] ;
  assign n28080 = ~n261 ;
  assign n7095 = n28080 & n7094 ;
  assign n16063 = x[64] & n7095 ;
  assign n17034 = n16063 & n28059 ;
  assign n28081 = ~n16063 ;
  assign n17035 = n28081 & n17033 ;
  assign n17036 = n17034 | n17035 ;
  assign n8767 = n6494 & n8706 ;
  assign n8705 = x[65] & n8645 ;
  assign n9901 = x[66] & n9278 ;
  assign n17037 = n8705 | n9901 ;
  assign n17038 = x[67] & n8643 ;
  assign n17039 = n17037 | n17038 ;
  assign n17040 = n8767 | n17039 ;
  assign n28082 = ~n17040 ;
  assign n17041 = x[17] & n28082 ;
  assign n17042 = n28039 & n17040 ;
  assign n17043 = n17041 | n17042 ;
  assign n17044 = n17036 | n17043 ;
  assign n17046 = n17036 & n17043 ;
  assign n28083 = ~n17046 ;
  assign n18068 = n17044 & n28083 ;
  assign n28084 = ~n18067 ;
  assign n18130 = n28084 & n18068 ;
  assign n28085 = ~n18068 ;
  assign n18131 = n18067 & n28085 ;
  assign n18132 = n18130 | n18131 ;
  assign n19081 = n18125 & n19080 ;
  assign n19082 = n18078 | n19081 ;
  assign n28086 = ~n18132 ;
  assign n19083 = n28086 & n19082 ;
  assign n28087 = ~n19082 ;
  assign n19306 = n18132 & n28087 ;
  assign n19307 = n19083 | n19306 ;
  assign n12710 = n3733 & n12695 ;
  assign n12663 = x[71] & n12633 ;
  assign n14405 = x[72] & n13533 ;
  assign n19308 = n12663 | n14405 ;
  assign n19309 = x[73] & n12631 ;
  assign n19310 = n19308 | n19309 ;
  assign n19311 = n12710 | n19310 ;
  assign n28088 = ~n19311 ;
  assign n19312 = x[11] & n28088 ;
  assign n19313 = n27892 & n19311 ;
  assign n19314 = n19312 | n19313 ;
  assign n19315 = n19307 & n19314 ;
  assign n19420 = n19307 | n19314 ;
  assign n28089 = ~n19315 ;
  assign n19421 = n28089 & n19420 ;
  assign n19409 = n19343 & n19407 ;
  assign n20351 = n19343 | n19407 ;
  assign n28090 = ~n19409 ;
  assign n20352 = n28090 & n20351 ;
  assign n20353 = n20349 & n20352 ;
  assign n20354 = n19346 | n20353 ;
  assign n20355 = n19414 & n20354 ;
  assign n20356 = n19336 | n20355 ;
  assign n20358 = n20356 & n20357 ;
  assign n20360 = n19326 | n20358 ;
  assign n28091 = ~n20360 ;
  assign n20361 = n19421 & n28091 ;
  assign n28092 = ~n19421 ;
  assign n20624 = n28092 & n20360 ;
  assign n20625 = n20361 | n20624 ;
  assign n20626 = n20623 & n20625 ;
  assign n20778 = n20623 | n20625 ;
  assign n28093 = ~n20626 ;
  assign n21182 = n28093 & n20778 ;
  assign n28094 = ~n20777 ;
  assign n21184 = n28094 & n21182 ;
  assign n28095 = ~n21182 ;
  assign n21668 = n20777 & n28095 ;
  assign n21669 = n21184 | n21668 ;
  assign n21670 = n21667 & n21669 ;
  assign n21870 = n21667 | n21669 ;
  assign n28096 = ~n21670 ;
  assign n21871 = n28096 & n21870 ;
  assign n22174 = n21855 & n22172 ;
  assign n22175 = n21713 | n22174 ;
  assign n21702 = n21697 | n21700 ;
  assign n22176 = n21702 & n28018 ;
  assign n22177 = n22175 & n22176 ;
  assign n22178 = n21703 | n22177 ;
  assign n22179 = n21863 & n22178 ;
  assign n22180 = n21690 | n22179 ;
  assign n22182 = n22180 & n22181 ;
  assign n22184 = n21680 | n22182 ;
  assign n28097 = ~n22184 ;
  assign n22185 = n21871 & n28097 ;
  assign n28098 = ~n21871 ;
  assign n22650 = n28098 & n22184 ;
  assign n22651 = n22185 | n22650 ;
  assign n507 = n505 & n506 ;
  assign n508 = n27644 | n507 ;
  assign n26634 = x[81] & x[82] ;
  assign n509 = x[81] | x[82] ;
  assign n28099 = ~n26634 ;
  assign n1000 = n28099 & n509 ;
  assign n1001 = n508 & n1000 ;
  assign n1002 = n508 | n1000 ;
  assign n28100 = ~n1001 ;
  assign n1003 = n28100 & n1002 ;
  assign n19665 = n1003 & n19656 ;
  assign n19774 = x[80] & n19723 ;
  assign n19846 = x[81] & n19829 ;
  assign n22652 = n19774 | n19846 ;
  assign n22653 = x[82] & n19655 ;
  assign n22654 = n22652 | n22653 ;
  assign n22655 = n19665 | n22654 ;
  assign n28101 = ~n22655 ;
  assign n22656 = x[2] & n28101 ;
  assign n22657 = n27790 & n22655 ;
  assign n22658 = n22656 | n22657 ;
  assign n28102 = ~n22658 ;
  assign n22659 = n22651 & n28102 ;
  assign n28103 = ~n22651 ;
  assign n22661 = n28103 & n22658 ;
  assign n22662 = n22659 | n22661 ;
  assign n22901 = n22673 | n22900 ;
  assign n22902 = n22662 & n22901 ;
  assign n27648 = n22662 | n22901 ;
  assign n28104 = ~n22902 ;
  assign n147 = n28104 & n27648 ;
  assign n18433 = n1270 & n18392 ;
  assign n18380 = x[78] & n18329 ;
  assign n18523 = x[79] & n18514 ;
  assign n21646 = n18380 | n18523 ;
  assign n21647 = x[80] & n18327 ;
  assign n21648 = n21646 | n21647 ;
  assign n21649 = n18433 | n21648 ;
  assign n28105 = ~n21649 ;
  assign n21650 = x[5] & n28105 ;
  assign n21651 = n27813 & n21649 ;
  assign n21652 = n21650 | n21651 ;
  assign n12698 = n2722 & n12695 ;
  assign n12636 = x[72] & n12633 ;
  assign n14406 = x[73] & n13533 ;
  assign n19292 = n12636 | n14406 ;
  assign n19293 = x[74] & n12631 ;
  assign n19294 = n19292 | n19293 ;
  assign n19295 = n12698 | n19294 ;
  assign n28106 = ~n19295 ;
  assign n19296 = x[11] & n28106 ;
  assign n19297 = n27892 & n19295 ;
  assign n19298 = n19296 | n19297 ;
  assign n18069 = n18067 & n18068 ;
  assign n18133 = n18128 & n18132 ;
  assign n18134 = n18069 | n18133 ;
  assign n10543 = n4790 & n10542 ;
  assign n10486 = x[69] & n10481 ;
  assign n11926 = x[70] & n11232 ;
  assign n18051 = n10486 | n11926 ;
  assign n18052 = x[71] & n10479 ;
  assign n18053 = n18051 | n18052 ;
  assign n18054 = n10543 | n18053 ;
  assign n28107 = ~n18054 ;
  assign n18055 = x[14] & n28107 ;
  assign n18056 = n27956 & n18054 ;
  assign n18057 = n18055 | n18056 ;
  assign n17045 = n16063 & n17033 ;
  assign n17047 = n17045 | n17046 ;
  assign n8768 = n6408 & n8706 ;
  assign n8685 = x[66] & n8645 ;
  assign n9853 = x[67] & n9278 ;
  assign n17048 = n8685 | n9853 ;
  assign n17049 = x[68] & n8643 ;
  assign n17050 = n17048 | n17049 ;
  assign n17051 = n8768 | n17050 ;
  assign n28108 = ~n17051 ;
  assign n17052 = x[17] & n28108 ;
  assign n17053 = n28039 & n17051 ;
  assign n17054 = n17052 | n17053 ;
  assign n16064 = x[20] & n28081 ;
  assign n262 = x[19] & x[20] ;
  assign n7096 = x[19] | x[20] ;
  assign n28109 = ~n262 ;
  assign n7097 = n28109 & n7096 ;
  assign n7162 = n7095 & n7097 ;
  assign n7222 = n6437 & n7162 ;
  assign n260 = x[18] & x[19] ;
  assign n7092 = x[18] | x[19] ;
  assign n28110 = ~n260 ;
  assign n7093 = n28110 & n7092 ;
  assign n28111 = ~n7095 ;
  assign n7647 = n7093 & n28111 ;
  assign n16065 = x[64] & n7647 ;
  assign n28112 = ~n7097 ;
  assign n7098 = n7095 & n28112 ;
  assign n16066 = x[65] & n7098 ;
  assign n16067 = n16065 | n16066 ;
  assign n16068 = n7222 | n16067 ;
  assign n28113 = ~n16068 ;
  assign n16069 = x[20] & n28113 ;
  assign n28114 = ~x[20] ;
  assign n16070 = n28114 & n16068 ;
  assign n16071 = n16069 | n16070 ;
  assign n28115 = ~n16071 ;
  assign n16072 = n16064 & n28115 ;
  assign n28116 = ~n16064 ;
  assign n17055 = n28116 & n16071 ;
  assign n17056 = n16072 | n17055 ;
  assign n28117 = ~n17054 ;
  assign n17057 = n28117 & n17056 ;
  assign n28118 = ~n17056 ;
  assign n17058 = n17054 & n28118 ;
  assign n17059 = n17057 | n17058 ;
  assign n28119 = ~n17059 ;
  assign n17061 = n17047 & n28119 ;
  assign n28120 = ~n17047 ;
  assign n18058 = n28120 & n17059 ;
  assign n18059 = n17061 | n18058 ;
  assign n18060 = n18057 & n18059 ;
  assign n18135 = n18057 | n18059 ;
  assign n28121 = ~n18060 ;
  assign n18136 = n28121 & n18135 ;
  assign n18137 = n18134 & n18136 ;
  assign n19301 = n18134 | n18136 ;
  assign n28122 = ~n18137 ;
  assign n19302 = n28122 & n19301 ;
  assign n28123 = ~n19298 ;
  assign n19303 = n28123 & n19302 ;
  assign n28124 = ~n19302 ;
  assign n19304 = n19298 & n28124 ;
  assign n19305 = n19303 | n19304 ;
  assign n19418 = n19325 & n19417 ;
  assign n19419 = n19326 | n19418 ;
  assign n19422 = n19419 & n19421 ;
  assign n19423 = n19315 | n19422 ;
  assign n19424 = n19305 | n19423 ;
  assign n19425 = n19305 & n19423 ;
  assign n28125 = ~n19425 ;
  assign n20602 = n19424 & n28125 ;
  assign n15313 = n1775 & n15308 ;
  assign n15250 = x[75] & n15246 ;
  assign n17310 = x[76] & n16288 ;
  assign n20603 = n15250 | n17310 ;
  assign n20604 = x[77] & n15244 ;
  assign n20605 = n20603 | n20604 ;
  assign n20606 = n15313 | n20605 ;
  assign n28126 = ~n20606 ;
  assign n20607 = x[8] & n28126 ;
  assign n20608 = n27845 & n20606 ;
  assign n20609 = n20607 | n20608 ;
  assign n28127 = ~n20609 ;
  assign n20610 = n20602 & n28127 ;
  assign n28128 = ~n20602 ;
  assign n21146 = n28128 & n20609 ;
  assign n21147 = n20610 | n21146 ;
  assign n21180 = n20774 & n21178 ;
  assign n21181 = n20636 | n21180 ;
  assign n21183 = n21181 & n21182 ;
  assign n21185 = n20626 | n21183 ;
  assign n21187 = n21147 | n21185 ;
  assign n21188 = n21147 & n21185 ;
  assign n28129 = ~n21188 ;
  assign n21656 = n21187 & n28129 ;
  assign n28130 = ~n21652 ;
  assign n21657 = n28130 & n21656 ;
  assign n28131 = ~n21656 ;
  assign n21659 = n21652 & n28131 ;
  assign n21660 = n21657 | n21659 ;
  assign n21868 = n21866 & n21867 ;
  assign n21869 = n21680 | n21868 ;
  assign n21872 = n21869 & n21871 ;
  assign n21873 = n21670 | n21872 ;
  assign n21874 = n21660 | n21873 ;
  assign n21875 = n21660 & n21873 ;
  assign n28132 = ~n21875 ;
  assign n22638 = n21874 & n28132 ;
  assign n510 = n508 & n509 ;
  assign n511 = n26634 | n510 ;
  assign n27639 = x[82] & x[83] ;
  assign n512 = x[82] | x[83] ;
  assign n28133 = ~n27639 ;
  assign n1054 = n28133 & n512 ;
  assign n28134 = ~n511 ;
  assign n1055 = n28134 & n1054 ;
  assign n28135 = ~n1054 ;
  assign n1056 = n511 & n28135 ;
  assign n1057 = n1055 | n1056 ;
  assign n19687 = n1057 & n19656 ;
  assign n19731 = x[81] & n19723 ;
  assign n19843 = x[82] & n19829 ;
  assign n22639 = n19731 | n19843 ;
  assign n22640 = x[83] & n19655 ;
  assign n22641 = n22639 | n22640 ;
  assign n22642 = n19687 | n22641 ;
  assign n28136 = ~n22642 ;
  assign n22643 = x[2] & n28136 ;
  assign n22644 = n27790 & n22642 ;
  assign n22645 = n22643 | n22644 ;
  assign n28137 = ~n22645 ;
  assign n22646 = n22638 & n28137 ;
  assign n28138 = ~n22638 ;
  assign n22648 = n28138 & n22645 ;
  assign n22649 = n22646 | n22648 ;
  assign n22660 = n22651 & n22658 ;
  assign n22903 = n22660 | n22902 ;
  assign n22904 = n22649 | n22903 ;
  assign n22905 = n22649 & n22903 ;
  assign n28139 = ~n22905 ;
  assign n148 = n22904 & n28139 ;
  assign n19084 = n18067 | n18068 ;
  assign n28140 = ~n18069 ;
  assign n19085 = n28140 & n19084 ;
  assign n19086 = n19082 & n19085 ;
  assign n19087 = n18069 | n19086 ;
  assign n28141 = ~n19087 ;
  assign n19088 = n18136 & n28141 ;
  assign n28142 = ~n18136 ;
  assign n19290 = n28142 & n19087 ;
  assign n19291 = n19088 | n19290 ;
  assign n19299 = n19291 | n19298 ;
  assign n19300 = n19291 & n19298 ;
  assign n28143 = ~n19300 ;
  assign n20338 = n19299 & n28143 ;
  assign n28144 = ~n19423 ;
  assign n20339 = n28144 & n20338 ;
  assign n28145 = ~n20338 ;
  assign n20612 = n19423 & n28145 ;
  assign n20613 = n20339 | n20612 ;
  assign n20614 = n20609 | n20613 ;
  assign n20615 = n20609 & n20613 ;
  assign n28146 = ~n20615 ;
  assign n20616 = n20614 & n28146 ;
  assign n28147 = ~n21185 ;
  assign n21186 = n20616 & n28147 ;
  assign n28148 = ~n20616 ;
  assign n21653 = n28148 & n21185 ;
  assign n21654 = n21186 | n21653 ;
  assign n21655 = n21652 & n21654 ;
  assign n21876 = n21655 | n21875 ;
  assign n18420 = n1029 & n18392 ;
  assign n18332 = x[79] & n18329 ;
  assign n18516 = x[80] & n18514 ;
  assign n21636 = n18332 | n18516 ;
  assign n21637 = x[81] & n18327 ;
  assign n21638 = n21636 | n21637 ;
  assign n21639 = n18420 | n21638 ;
  assign n28149 = ~n21639 ;
  assign n21640 = x[5] & n28149 ;
  assign n21641 = n27813 & n21639 ;
  assign n21642 = n21640 | n21641 ;
  assign n15342 = n2084 & n15308 ;
  assign n15251 = x[76] & n15246 ;
  assign n17280 = x[77] & n16288 ;
  assign n20589 = n15251 | n17280 ;
  assign n20590 = x[78] & n15244 ;
  assign n20591 = n20589 | n20590 ;
  assign n20592 = n15342 | n20591 ;
  assign n28150 = ~n20592 ;
  assign n20593 = x[8] & n28150 ;
  assign n20594 = n27845 & n20592 ;
  assign n20595 = n20593 | n20594 ;
  assign n19426 = n19300 | n19425 ;
  assign n12699 = n3289 & n12695 ;
  assign n12650 = x[73] & n12633 ;
  assign n14356 = x[74] & n13533 ;
  assign n19280 = n12650 | n14356 ;
  assign n19281 = x[75] & n12631 ;
  assign n19282 = n19280 | n19281 ;
  assign n19283 = n12699 | n19282 ;
  assign n28151 = ~n19283 ;
  assign n19284 = x[11] & n28151 ;
  assign n19285 = n27892 & n19283 ;
  assign n19286 = n19284 | n19285 ;
  assign n18138 = n18060 | n18137 ;
  assign n17060 = n17047 & n17059 ;
  assign n17062 = n17054 & n17056 ;
  assign n17063 = n17060 | n17062 ;
  assign n16073 = n16064 & n16071 ;
  assign n7223 = n6466 & n7162 ;
  assign n7099 = n28111 & n7097 ;
  assign n28152 = ~n7093 ;
  assign n7100 = n28152 & n7099 ;
  assign n7159 = x[64] & n7100 ;
  assign n7728 = x[65] & n7647 ;
  assign n16074 = n7159 | n7728 ;
  assign n16075 = x[66] & n7098 ;
  assign n16076 = n16074 | n16075 ;
  assign n16077 = n7223 | n16076 ;
  assign n28153 = ~n16077 ;
  assign n16078 = x[20] & n28153 ;
  assign n16079 = n28114 & n16077 ;
  assign n16080 = n16078 | n16079 ;
  assign n16081 = n16073 | n16080 ;
  assign n16082 = n16073 & n16080 ;
  assign n28154 = ~n16082 ;
  assign n17005 = n16081 & n28154 ;
  assign n8723 = n6379 & n8706 ;
  assign n8647 = x[67] & n8645 ;
  assign n9895 = x[68] & n9278 ;
  assign n17006 = n8647 | n9895 ;
  assign n17007 = x[69] & n8643 ;
  assign n17008 = n17006 | n17007 ;
  assign n17009 = n8723 | n17008 ;
  assign n28155 = ~n17009 ;
  assign n17010 = x[17] & n28155 ;
  assign n17011 = n28039 & n17009 ;
  assign n17012 = n17010 | n17011 ;
  assign n17013 = n17005 & n17012 ;
  assign n17064 = n17005 | n17012 ;
  assign n28156 = ~n17013 ;
  assign n18038 = n28156 & n17064 ;
  assign n28157 = ~n18038 ;
  assign n18039 = n17063 & n28157 ;
  assign n17065 = n17063 & n17064 ;
  assign n17066 = n17013 | n17065 ;
  assign n28158 = ~n17066 ;
  assign n18040 = n17064 & n28158 ;
  assign n18041 = n18039 | n18040 ;
  assign n10545 = n3701 & n10542 ;
  assign n10514 = x[70] & n10481 ;
  assign n11921 = x[71] & n11232 ;
  assign n18042 = n10514 | n11921 ;
  assign n18043 = x[72] & n10479 ;
  assign n18044 = n18042 | n18043 ;
  assign n18045 = n10545 | n18044 ;
  assign n28159 = ~n18045 ;
  assign n18046 = x[14] & n28159 ;
  assign n18047 = n27956 & n18045 ;
  assign n18048 = n18046 | n18047 ;
  assign n28160 = ~n18048 ;
  assign n18049 = n18041 & n28160 ;
  assign n28161 = ~n18041 ;
  assign n19091 = n28161 & n18048 ;
  assign n19092 = n18049 | n19091 ;
  assign n28162 = ~n18138 ;
  assign n19094 = n28162 & n19092 ;
  assign n28163 = ~n19092 ;
  assign n19287 = n18138 & n28163 ;
  assign n19288 = n19094 | n19287 ;
  assign n19289 = n19286 & n19288 ;
  assign n19427 = n19286 | n19288 ;
  assign n28164 = ~n19289 ;
  assign n19428 = n28164 & n19427 ;
  assign n19429 = n19426 & n19428 ;
  assign n20596 = n19426 | n19428 ;
  assign n28165 = ~n19429 ;
  assign n20597 = n28165 & n20596 ;
  assign n28166 = ~n20595 ;
  assign n20599 = n28166 & n20597 ;
  assign n28167 = ~n20597 ;
  assign n20600 = n20595 & n28167 ;
  assign n20601 = n20599 | n20600 ;
  assign n20611 = n20602 & n20609 ;
  assign n20779 = n20777 & n20778 ;
  assign n20780 = n20626 | n20779 ;
  assign n20781 = n20616 & n20780 ;
  assign n20782 = n20611 | n20781 ;
  assign n20783 = n20601 | n20782 ;
  assign n20784 = n20601 & n20782 ;
  assign n28168 = ~n20784 ;
  assign n21877 = n20783 & n28168 ;
  assign n28169 = ~n21642 ;
  assign n21879 = n28169 & n21877 ;
  assign n28170 = ~n21877 ;
  assign n22190 = n21642 & n28170 ;
  assign n22191 = n21879 | n22190 ;
  assign n28171 = ~n22191 ;
  assign n22192 = n21876 & n28171 ;
  assign n28172 = ~n21876 ;
  assign n22625 = n28172 & n22191 ;
  assign n22626 = n22192 | n22625 ;
  assign n513 = n511 & n512 ;
  assign n514 = n27639 | n513 ;
  assign n26534 = x[83] & x[84] ;
  assign n515 = x[83] | x[84] ;
  assign n28173 = ~n26534 ;
  assign n1290 = n28173 & n515 ;
  assign n1291 = n514 & n1290 ;
  assign n1292 = n514 | n1290 ;
  assign n28174 = ~n1291 ;
  assign n1293 = n28174 & n1292 ;
  assign n19669 = n1293 & n19656 ;
  assign n19748 = x[82] & n19723 ;
  assign n19889 = x[83] & n19829 ;
  assign n22627 = n19748 | n19889 ;
  assign n22628 = x[84] & n19655 ;
  assign n22629 = n22627 | n22628 ;
  assign n22630 = n19669 | n22629 ;
  assign n28175 = ~n22630 ;
  assign n22631 = x[2] & n28175 ;
  assign n22632 = n27790 & n22630 ;
  assign n22633 = n22631 | n22632 ;
  assign n28176 = ~n22633 ;
  assign n22634 = n22626 & n28176 ;
  assign n28177 = ~n22626 ;
  assign n22636 = n28177 & n22633 ;
  assign n22637 = n22634 | n22636 ;
  assign n22647 = n22638 & n22645 ;
  assign n22906 = n22647 | n22905 ;
  assign n22907 = n22637 & n22906 ;
  assign n27651 = n22637 | n22906 ;
  assign n28178 = ~n22907 ;
  assign n149 = n28178 & n27651 ;
  assign n20598 = n20595 & n20597 ;
  assign n20785 = n20598 | n20784 ;
  assign n15316 = n1741 & n15308 ;
  assign n15252 = x[77] & n15246 ;
  assign n17330 = x[78] & n16288 ;
  assign n20579 = n15252 | n17330 ;
  assign n20580 = x[79] & n15244 ;
  assign n20581 = n20579 | n20580 ;
  assign n20582 = n15316 | n20581 ;
  assign n28179 = ~n20582 ;
  assign n20583 = x[8] & n28179 ;
  assign n20584 = n27845 & n20582 ;
  assign n20585 = n20583 | n20584 ;
  assign n19430 = n19289 | n19429 ;
  assign n12725 = n2750 & n12695 ;
  assign n12643 = x[74] & n12633 ;
  assign n14368 = x[75] & n13533 ;
  assign n19270 = n12643 | n14368 ;
  assign n19271 = x[76] & n12631 ;
  assign n19272 = n19270 | n19271 ;
  assign n19273 = n12725 | n19272 ;
  assign n28180 = ~n19273 ;
  assign n19274 = x[11] & n28180 ;
  assign n19275 = n27892 & n19273 ;
  assign n19276 = n19274 | n19275 ;
  assign n8707 = n5976 & n8706 ;
  assign n8667 = x[68] & n8645 ;
  assign n9900 = x[69] & n9278 ;
  assign n16995 = n8667 | n9900 ;
  assign n16996 = x[70] & n8643 ;
  assign n16997 = n16995 | n16996 ;
  assign n16998 = n8707 | n16997 ;
  assign n16999 = x[17] | n16998 ;
  assign n17000 = x[17] & n16998 ;
  assign n28181 = ~n17000 ;
  assign n17001 = n16999 & n28181 ;
  assign n27773 = x[20] & x[21] ;
  assign n5234 = x[20] | x[21] ;
  assign n28182 = ~n27773 ;
  assign n5235 = n28182 & n5234 ;
  assign n15005 = x[64] & n5235 ;
  assign n16083 = n15005 & n28154 ;
  assign n28183 = ~n15005 ;
  assign n16084 = n28183 & n16082 ;
  assign n16085 = n16083 | n16084 ;
  assign n7224 = n6494 & n7162 ;
  assign n7160 = x[65] & n7100 ;
  assign n7671 = x[66] & n7647 ;
  assign n16086 = n7160 | n7671 ;
  assign n16087 = x[67] & n7098 ;
  assign n16088 = n16086 | n16087 ;
  assign n16089 = n7224 | n16088 ;
  assign n28184 = ~n16089 ;
  assign n16090 = x[20] & n28184 ;
  assign n16091 = n28114 & n16089 ;
  assign n16092 = n16090 | n16091 ;
  assign n28185 = ~n16092 ;
  assign n16093 = n16085 & n28185 ;
  assign n28186 = ~n16085 ;
  assign n17002 = n28186 & n16092 ;
  assign n17003 = n16093 | n17002 ;
  assign n17004 = n17001 & n17003 ;
  assign n17067 = n17001 | n17003 ;
  assign n28187 = ~n17004 ;
  assign n17068 = n28187 & n17067 ;
  assign n17069 = n17066 & n17068 ;
  assign n18028 = n17066 | n17068 ;
  assign n28188 = ~n17069 ;
  assign n18029 = n28188 & n18028 ;
  assign n10547 = n3733 & n10542 ;
  assign n10488 = x[71] & n10481 ;
  assign n11925 = x[72] & n11232 ;
  assign n18030 = n10488 | n11925 ;
  assign n18031 = x[73] & n10479 ;
  assign n18032 = n18030 | n18031 ;
  assign n18033 = n10547 | n18032 ;
  assign n28189 = ~n18033 ;
  assign n18034 = x[14] & n28189 ;
  assign n18035 = n27956 & n18033 ;
  assign n18036 = n18034 | n18035 ;
  assign n18037 = n18029 & n18036 ;
  assign n18142 = n18029 | n18036 ;
  assign n28190 = ~n18037 ;
  assign n18143 = n28190 & n18142 ;
  assign n18050 = n18041 & n18048 ;
  assign n19089 = n18135 & n19087 ;
  assign n19090 = n18060 | n19089 ;
  assign n19093 = n19090 & n19092 ;
  assign n19095 = n18050 | n19093 ;
  assign n28191 = ~n19095 ;
  assign n19096 = n18143 & n28191 ;
  assign n28192 = ~n18143 ;
  assign n19277 = n28192 & n19095 ;
  assign n19278 = n19096 | n19277 ;
  assign n19279 = n19276 & n19278 ;
  assign n19431 = n19276 | n19278 ;
  assign n28193 = ~n19279 ;
  assign n20368 = n28193 & n19431 ;
  assign n28194 = ~n19430 ;
  assign n20370 = n28194 & n20368 ;
  assign n28195 = ~n20368 ;
  assign n20586 = n19430 & n28195 ;
  assign n20587 = n20370 | n20586 ;
  assign n20588 = n20585 & n20587 ;
  assign n20786 = n20585 | n20587 ;
  assign n28196 = ~n20588 ;
  assign n20787 = n28196 & n20786 ;
  assign n20788 = n20785 & n20787 ;
  assign n21622 = n20785 | n20787 ;
  assign n28197 = ~n20788 ;
  assign n21623 = n28197 & n21622 ;
  assign n18403 = n1003 & n18392 ;
  assign n18363 = x[80] & n18329 ;
  assign n18558 = x[81] & n18514 ;
  assign n21624 = n18363 | n18558 ;
  assign n21625 = x[82] & n18327 ;
  assign n21626 = n21624 | n21625 ;
  assign n21627 = n18403 | n21626 ;
  assign n28198 = ~n21627 ;
  assign n21628 = x[5] & n28198 ;
  assign n21629 = n27813 & n21627 ;
  assign n21630 = n21628 | n21629 ;
  assign n28199 = ~n21630 ;
  assign n21633 = n21623 & n28199 ;
  assign n28200 = ~n21623 ;
  assign n21634 = n28200 & n21630 ;
  assign n21635 = n21633 | n21634 ;
  assign n21143 = n20595 | n20597 ;
  assign n28201 = ~n20598 ;
  assign n21144 = n28201 & n21143 ;
  assign n28202 = ~n20782 ;
  assign n21145 = n28202 & n21144 ;
  assign n28203 = ~n21144 ;
  assign n21643 = n20782 & n28203 ;
  assign n21644 = n21145 | n21643 ;
  assign n21645 = n21642 & n21644 ;
  assign n21878 = n21642 & n21877 ;
  assign n21880 = n21642 | n21877 ;
  assign n28204 = ~n21878 ;
  assign n21881 = n28204 & n21880 ;
  assign n21882 = n21876 & n21881 ;
  assign n21883 = n21645 | n21882 ;
  assign n21884 = n21635 | n21883 ;
  assign n21885 = n21635 & n21883 ;
  assign n28205 = ~n21885 ;
  assign n22613 = n21884 & n28205 ;
  assign n516 = n514 & n515 ;
  assign n517 = n26534 | n516 ;
  assign n27637 = x[84] & x[85] ;
  assign n518 = x[84] | x[85] ;
  assign n28206 = ~n27637 ;
  assign n1236 = n28206 & n518 ;
  assign n1237 = n517 | n1236 ;
  assign n1238 = n517 & n1236 ;
  assign n28207 = ~n1238 ;
  assign n1239 = n1237 & n28207 ;
  assign n19670 = n1239 & n19656 ;
  assign n19742 = x[83] & n19723 ;
  assign n19844 = x[84] & n19829 ;
  assign n22614 = n19742 | n19844 ;
  assign n22615 = x[85] & n19655 ;
  assign n22616 = n22614 | n22615 ;
  assign n22617 = n19670 | n22616 ;
  assign n28208 = ~n22617 ;
  assign n22618 = x[2] & n28208 ;
  assign n22619 = n27790 & n22617 ;
  assign n22620 = n22618 | n22619 ;
  assign n28209 = ~n22620 ;
  assign n22621 = n22613 & n28209 ;
  assign n28210 = ~n22613 ;
  assign n22623 = n28210 & n22620 ;
  assign n22624 = n22621 | n22623 ;
  assign n22635 = n22626 & n22633 ;
  assign n22908 = n22635 | n22907 ;
  assign n22909 = n22624 | n22908 ;
  assign n22910 = n22624 & n22908 ;
  assign n28211 = ~n22910 ;
  assign n150 = n22909 & n28211 ;
  assign n22622 = n22613 & n22620 ;
  assign n22911 = n22622 | n22910 ;
  assign n20789 = n20588 | n20788 ;
  assign n15318 = n1270 & n15308 ;
  assign n15268 = x[78] & n15246 ;
  assign n17282 = x[79] & n16288 ;
  assign n20569 = n15268 | n17282 ;
  assign n20570 = x[80] & n15244 ;
  assign n20571 = n20569 | n20570 ;
  assign n20572 = n15318 | n20571 ;
  assign n28212 = ~n20572 ;
  assign n20573 = x[8] & n28212 ;
  assign n20574 = n27845 & n20572 ;
  assign n20575 = n20573 | n20574 ;
  assign n12731 = n1775 & n12695 ;
  assign n12658 = x[75] & n12633 ;
  assign n14397 = x[76] & n13533 ;
  assign n19262 = n12658 | n14397 ;
  assign n19263 = x[77] & n12631 ;
  assign n19264 = n19262 | n19263 ;
  assign n19265 = n12731 | n19264 ;
  assign n28213 = ~n19265 ;
  assign n19266 = x[11] & n28213 ;
  assign n19267 = n27892 & n19265 ;
  assign n19268 = n19266 | n19267 ;
  assign n18139 = n18041 | n18048 ;
  assign n18140 = n18138 & n18139 ;
  assign n18141 = n18050 | n18140 ;
  assign n18144 = n18141 & n18143 ;
  assign n18145 = n18037 | n18144 ;
  assign n17070 = n17004 | n17069 ;
  assign n8708 = n4790 & n8706 ;
  assign n8671 = x[69] & n8645 ;
  assign n9882 = x[70] & n9278 ;
  assign n16985 = n8671 | n9882 ;
  assign n16986 = x[71] & n8643 ;
  assign n16987 = n16985 | n16986 ;
  assign n16988 = n8708 | n16987 ;
  assign n16989 = x[17] | n16988 ;
  assign n16990 = x[17] & n16988 ;
  assign n28214 = ~n16990 ;
  assign n16991 = n16989 & n28214 ;
  assign n16094 = n16085 & n16092 ;
  assign n16095 = n15005 & n16082 ;
  assign n16096 = n16094 | n16095 ;
  assign n7225 = n6408 & n7162 ;
  assign n7161 = x[66] & n7100 ;
  assign n7730 = x[67] & n7647 ;
  assign n16097 = n7161 | n7730 ;
  assign n16098 = x[68] & n7098 ;
  assign n16099 = n16097 | n16098 ;
  assign n16100 = n7225 | n16099 ;
  assign n28215 = ~n16100 ;
  assign n16101 = x[20] & n28215 ;
  assign n16102 = n28114 & n16100 ;
  assign n16103 = n16101 | n16102 ;
  assign n15006 = x[23] & n28183 ;
  assign n27774 = x[22] & x[23] ;
  assign n5236 = x[22] | x[23] ;
  assign n28216 = ~n27774 ;
  assign n5237 = n28216 & n5236 ;
  assign n5302 = n5235 & n5237 ;
  assign n6451 = n5302 & n6437 ;
  assign n27770 = x[21] & x[22] ;
  assign n5232 = x[21] | x[22] ;
  assign n28217 = ~n27770 ;
  assign n5233 = n28217 & n5232 ;
  assign n28218 = ~n5235 ;
  assign n6179 = n5233 & n28218 ;
  assign n15007 = x[64] & n6179 ;
  assign n28219 = ~n5237 ;
  assign n5238 = n5235 & n28219 ;
  assign n15008 = x[65] & n5238 ;
  assign n15009 = n15007 | n15008 ;
  assign n15010 = n6451 | n15009 ;
  assign n28220 = ~n15010 ;
  assign n15011 = x[23] & n28220 ;
  assign n28221 = ~x[23] ;
  assign n15012 = n28221 & n15010 ;
  assign n15013 = n15011 | n15012 ;
  assign n28222 = ~n15013 ;
  assign n15014 = n15006 & n28222 ;
  assign n28223 = ~n15006 ;
  assign n16104 = n28223 & n15013 ;
  assign n16105 = n15014 | n16104 ;
  assign n28224 = ~n16103 ;
  assign n16106 = n28224 & n16105 ;
  assign n28225 = ~n16105 ;
  assign n16107 = n16103 & n28225 ;
  assign n16108 = n16106 | n16107 ;
  assign n16109 = n16096 & n16108 ;
  assign n16992 = n16096 | n16108 ;
  assign n28226 = ~n16109 ;
  assign n16993 = n28226 & n16992 ;
  assign n16994 = n16991 & n16993 ;
  assign n17071 = n16991 | n16993 ;
  assign n28227 = ~n16994 ;
  assign n17072 = n28227 & n17071 ;
  assign n28228 = ~n17070 ;
  assign n17073 = n28228 & n17072 ;
  assign n28229 = ~n17072 ;
  assign n18014 = n17070 & n28229 ;
  assign n18015 = n17073 | n18014 ;
  assign n10561 = n2722 & n10542 ;
  assign n10511 = x[72] & n10481 ;
  assign n11900 = x[73] & n11232 ;
  assign n18016 = n10511 | n11900 ;
  assign n18017 = x[74] & n10479 ;
  assign n18018 = n18016 | n18017 ;
  assign n18019 = n10561 | n18018 ;
  assign n28230 = ~n18019 ;
  assign n18020 = x[14] & n28230 ;
  assign n18021 = n27956 & n18019 ;
  assign n18022 = n18020 | n18021 ;
  assign n18023 = n18015 | n18022 ;
  assign n18024 = n18015 & n18022 ;
  assign n28231 = ~n18024 ;
  assign n19071 = n18023 & n28231 ;
  assign n28232 = ~n18145 ;
  assign n19072 = n28232 & n19071 ;
  assign n28233 = ~n19071 ;
  assign n19434 = n18145 & n28233 ;
  assign n19435 = n19072 | n19434 ;
  assign n19436 = n19268 & n19435 ;
  assign n28234 = ~n18022 ;
  assign n18025 = n18015 & n28234 ;
  assign n28235 = ~n18015 ;
  assign n18026 = n28235 & n18022 ;
  assign n18027 = n18025 | n18026 ;
  assign n18146 = n18027 | n18145 ;
  assign n18147 = n18027 & n18145 ;
  assign n28236 = ~n18147 ;
  assign n19261 = n18146 & n28236 ;
  assign n19437 = n19261 | n19268 ;
  assign n28237 = ~n19436 ;
  assign n19438 = n28237 & n19437 ;
  assign n20337 = n19298 & n19302 ;
  assign n20362 = n19420 & n20360 ;
  assign n20363 = n19315 | n20362 ;
  assign n20364 = n20338 & n20363 ;
  assign n20365 = n20337 | n20364 ;
  assign n20366 = n19427 & n20365 ;
  assign n20367 = n19289 | n20366 ;
  assign n20369 = n20367 & n20368 ;
  assign n20371 = n19279 | n20369 ;
  assign n28238 = ~n20371 ;
  assign n20372 = n19438 & n28238 ;
  assign n28239 = ~n19438 ;
  assign n20576 = n28239 & n20371 ;
  assign n20577 = n20372 | n20576 ;
  assign n20578 = n20575 & n20577 ;
  assign n20790 = n20575 | n20577 ;
  assign n28240 = ~n20578 ;
  assign n21194 = n28240 & n20790 ;
  assign n28241 = ~n20789 ;
  assign n21196 = n28241 & n21194 ;
  assign n28242 = ~n21194 ;
  assign n21609 = n20789 & n28242 ;
  assign n21610 = n21196 | n21609 ;
  assign n18444 = n1057 & n18392 ;
  assign n18336 = x[81] & n18329 ;
  assign n18542 = x[82] & n18514 ;
  assign n21611 = n18336 | n18542 ;
  assign n21612 = x[83] & n18327 ;
  assign n21613 = n21611 | n21612 ;
  assign n21614 = n18444 | n21613 ;
  assign n28243 = ~n21614 ;
  assign n21615 = x[5] & n28243 ;
  assign n21616 = n27813 & n21614 ;
  assign n21617 = n21615 | n21616 ;
  assign n21619 = n21610 & n21617 ;
  assign n21620 = n21610 | n21617 ;
  assign n28244 = ~n21619 ;
  assign n21621 = n28244 & n21620 ;
  assign n21632 = n21623 & n21630 ;
  assign n21631 = n21623 | n21630 ;
  assign n28245 = ~n21632 ;
  assign n22128 = n21631 & n28245 ;
  assign n21658 = n21652 & n21656 ;
  assign n22129 = n21652 | n21656 ;
  assign n28246 = ~n21658 ;
  assign n22130 = n28246 & n22129 ;
  assign n22186 = n21870 & n22184 ;
  assign n22187 = n21670 | n22186 ;
  assign n22188 = n22130 & n22187 ;
  assign n22189 = n21655 | n22188 ;
  assign n22193 = n22189 & n22191 ;
  assign n22194 = n21645 | n22193 ;
  assign n22195 = n22128 & n22194 ;
  assign n22196 = n21632 | n22195 ;
  assign n28247 = ~n22196 ;
  assign n22197 = n21621 & n28247 ;
  assign n28248 = ~n21621 ;
  assign n22602 = n28248 & n22196 ;
  assign n22603 = n22197 | n22602 ;
  assign n519 = n517 & n518 ;
  assign n520 = n27637 | n519 ;
  assign n26427 = x[85] & x[86] ;
  assign n521 = x[85] | x[86] ;
  assign n28249 = ~n26427 ;
  assign n1210 = n28249 & n521 ;
  assign n1211 = n520 & n1210 ;
  assign n1212 = n520 | n1210 ;
  assign n28250 = ~n1211 ;
  assign n1213 = n28250 & n1212 ;
  assign n19672 = n1213 & n19656 ;
  assign n19733 = x[84] & n19723 ;
  assign n19852 = x[85] & n19829 ;
  assign n22604 = n19733 | n19852 ;
  assign n22605 = x[86] & n19655 ;
  assign n22606 = n22604 | n22605 ;
  assign n22607 = n19672 | n22606 ;
  assign n28251 = ~n22607 ;
  assign n22608 = x[2] & n28251 ;
  assign n22609 = n27790 & n22607 ;
  assign n22610 = n22608 | n22609 ;
  assign n22611 = n22603 | n22610 ;
  assign n22612 = n22603 & n22610 ;
  assign n28252 = ~n22612 ;
  assign n22912 = n22611 & n28252 ;
  assign n22913 = n22911 & n22912 ;
  assign n27654 = n22911 | n22912 ;
  assign n28253 = ~n22913 ;
  assign n151 = n28253 & n27654 ;
  assign n21189 = n20615 | n21188 ;
  assign n21190 = n21144 & n21189 ;
  assign n21191 = n20598 | n21190 ;
  assign n21192 = n20786 & n21191 ;
  assign n21193 = n20588 | n21192 ;
  assign n21195 = n21193 & n21194 ;
  assign n21197 = n20578 | n21195 ;
  assign n15367 = n1029 & n15308 ;
  assign n15282 = x[79] & n15246 ;
  assign n17287 = x[80] & n16288 ;
  assign n20559 = n15282 | n17287 ;
  assign n20560 = x[81] & n15244 ;
  assign n20561 = n20559 | n20560 ;
  assign n20562 = n15367 | n20561 ;
  assign n28254 = ~n20562 ;
  assign n20563 = x[8] & n28254 ;
  assign n20564 = n27845 & n20562 ;
  assign n20565 = n20563 | n20564 ;
  assign n12737 = n2084 & n12695 ;
  assign n12689 = x[76] & n12633 ;
  assign n14357 = x[77] & n13533 ;
  assign n19248 = n12689 | n14357 ;
  assign n19249 = x[78] & n12631 ;
  assign n19250 = n19248 | n19249 ;
  assign n19251 = n12737 | n19250 ;
  assign n28255 = ~n19251 ;
  assign n19252 = x[11] & n28255 ;
  assign n19253 = n27892 & n19251 ;
  assign n19254 = n19252 | n19253 ;
  assign n18148 = n18024 | n18147 ;
  assign n10548 = n3289 & n10542 ;
  assign n10538 = x[73] & n10481 ;
  assign n11911 = x[74] & n11232 ;
  assign n18004 = n10538 | n11911 ;
  assign n18005 = x[75] & n10479 ;
  assign n18006 = n18004 | n18005 ;
  assign n18007 = n10548 | n18006 ;
  assign n28256 = ~n18007 ;
  assign n18008 = x[14] & n28256 ;
  assign n18009 = n27956 & n18007 ;
  assign n18010 = n18008 | n18009 ;
  assign n17074 = n17070 & n17072 ;
  assign n17075 = n16994 | n17074 ;
  assign n16110 = n16103 & n16105 ;
  assign n16111 = n16109 | n16110 ;
  assign n15015 = n15006 & n15013 ;
  assign n6480 = n5302 & n6466 ;
  assign n5239 = n28218 & n5237 ;
  assign n28257 = ~n5233 ;
  assign n5240 = n28257 & n5239 ;
  assign n5256 = x[64] & n5240 ;
  assign n6230 = x[65] & n6179 ;
  assign n15016 = n5256 | n6230 ;
  assign n15017 = x[66] & n5238 ;
  assign n15018 = n15016 | n15017 ;
  assign n15019 = n6480 | n15018 ;
  assign n28258 = ~n15019 ;
  assign n15020 = x[23] & n28258 ;
  assign n15021 = n28221 & n15019 ;
  assign n15022 = n15020 | n15021 ;
  assign n15023 = n15015 | n15022 ;
  assign n15024 = n15015 & n15022 ;
  assign n28259 = ~n15024 ;
  assign n16054 = n15023 & n28259 ;
  assign n7220 = n6379 & n7162 ;
  assign n7126 = x[67] & n7100 ;
  assign n7707 = x[68] & n7647 ;
  assign n16055 = n7126 | n7707 ;
  assign n16056 = x[69] & n7098 ;
  assign n16057 = n16055 | n16056 ;
  assign n16058 = n7220 | n16057 ;
  assign n28260 = ~n16058 ;
  assign n16059 = x[20] & n28260 ;
  assign n16060 = n28114 & n16058 ;
  assign n16061 = n16059 | n16060 ;
  assign n16062 = n16054 & n16061 ;
  assign n16112 = n16054 | n16061 ;
  assign n28261 = ~n16062 ;
  assign n16972 = n28261 & n16112 ;
  assign n28262 = ~n16972 ;
  assign n16973 = n16111 & n28262 ;
  assign n16113 = n16111 & n16112 ;
  assign n16114 = n16062 | n16113 ;
  assign n28263 = ~n16114 ;
  assign n16974 = n16112 & n28263 ;
  assign n16975 = n16973 | n16974 ;
  assign n8716 = n3701 & n8706 ;
  assign n8648 = x[70] & n8645 ;
  assign n9899 = x[71] & n9278 ;
  assign n16976 = n8648 | n9899 ;
  assign n16977 = x[72] & n8643 ;
  assign n16978 = n16976 | n16977 ;
  assign n16979 = n8716 | n16978 ;
  assign n28264 = ~n16979 ;
  assign n16980 = x[17] & n28264 ;
  assign n16981 = n28039 & n16979 ;
  assign n16982 = n16980 | n16981 ;
  assign n28265 = ~n16982 ;
  assign n16983 = n16975 & n28265 ;
  assign n28266 = ~n16975 ;
  assign n17773 = n28266 & n16982 ;
  assign n17774 = n16983 | n17773 ;
  assign n17775 = n17075 & n17774 ;
  assign n18149 = n17075 | n17774 ;
  assign n28267 = ~n17775 ;
  assign n18150 = n28267 & n18149 ;
  assign n18151 = n18010 & n18150 ;
  assign n18152 = n18010 | n18150 ;
  assign n28268 = ~n18151 ;
  assign n18153 = n28268 & n18152 ;
  assign n18154 = n18148 & n18153 ;
  assign n19255 = n18148 | n18153 ;
  assign n28269 = ~n18154 ;
  assign n19256 = n28269 & n19255 ;
  assign n28270 = ~n19254 ;
  assign n19258 = n28270 & n19256 ;
  assign n28271 = ~n19256 ;
  assign n19259 = n19254 & n28271 ;
  assign n19260 = n19258 | n19259 ;
  assign n19269 = n19261 & n19268 ;
  assign n19432 = n19430 & n19431 ;
  assign n19433 = n19279 | n19432 ;
  assign n19439 = n19433 & n19438 ;
  assign n19440 = n19269 | n19439 ;
  assign n19441 = n19260 | n19440 ;
  assign n19442 = n19260 & n19440 ;
  assign n28272 = ~n19442 ;
  assign n20793 = n19441 & n28272 ;
  assign n28273 = ~n20565 ;
  assign n20795 = n28273 & n20793 ;
  assign n28274 = ~n20793 ;
  assign n21198 = n20565 & n28274 ;
  assign n21199 = n20795 | n21198 ;
  assign n21200 = n21197 | n21199 ;
  assign n21201 = n21197 & n21199 ;
  assign n28275 = ~n21201 ;
  assign n21596 = n21200 & n28275 ;
  assign n18396 = n1293 & n18392 ;
  assign n18337 = x[82] & n18329 ;
  assign n18524 = x[83] & n18514 ;
  assign n21597 = n18337 | n18524 ;
  assign n21598 = x[84] & n18327 ;
  assign n21599 = n21597 | n21598 ;
  assign n21600 = n18396 | n21599 ;
  assign n28276 = ~n21600 ;
  assign n21601 = x[5] & n28276 ;
  assign n21602 = n27813 & n21600 ;
  assign n21603 = n21601 | n21602 ;
  assign n28277 = ~n21603 ;
  assign n21606 = n21596 & n28277 ;
  assign n28278 = ~n21596 ;
  assign n21607 = n28278 & n21603 ;
  assign n21608 = n21606 | n21607 ;
  assign n21886 = n21632 | n21885 ;
  assign n21887 = n21621 & n21886 ;
  assign n21888 = n21619 | n21887 ;
  assign n21889 = n21608 | n21888 ;
  assign n21890 = n21608 & n21888 ;
  assign n28279 = ~n21890 ;
  assign n22590 = n21889 & n28279 ;
  assign n522 = n520 & n521 ;
  assign n523 = n26427 | n522 ;
  assign n27636 = x[86] & x[87] ;
  assign n524 = x[86] | x[87] ;
  assign n28280 = ~n27636 ;
  assign n1519 = n28280 & n524 ;
  assign n28281 = ~n523 ;
  assign n1520 = n28281 & n1519 ;
  assign n28282 = ~n1519 ;
  assign n1521 = n523 & n28282 ;
  assign n1522 = n1520 | n1521 ;
  assign n19696 = n1522 & n19656 ;
  assign n19738 = x[85] & n19723 ;
  assign n19848 = x[86] & n19829 ;
  assign n22591 = n19738 | n19848 ;
  assign n22592 = x[87] & n19655 ;
  assign n22593 = n22591 | n22592 ;
  assign n22594 = n19696 | n22593 ;
  assign n28283 = ~n22594 ;
  assign n22595 = x[2] & n28283 ;
  assign n22596 = n27790 & n22594 ;
  assign n22597 = n22595 | n22596 ;
  assign n28284 = ~n22597 ;
  assign n22598 = n22590 & n28284 ;
  assign n28285 = ~n22590 ;
  assign n22600 = n28285 & n22597 ;
  assign n22601 = n22598 | n22600 ;
  assign n22914 = n22612 | n22913 ;
  assign n22915 = n22601 | n22914 ;
  assign n22916 = n22601 & n22914 ;
  assign n28286 = ~n22916 ;
  assign n152 = n22915 & n28286 ;
  assign n21605 = n21596 & n21603 ;
  assign n21891 = n21605 | n21890 ;
  assign n18425 = n1239 & n18392 ;
  assign n18390 = x[83] & n18329 ;
  assign n18531 = x[84] & n18514 ;
  assign n21586 = n18390 | n18531 ;
  assign n21587 = x[85] & n18327 ;
  assign n21588 = n21586 | n21587 ;
  assign n21589 = n18425 | n21588 ;
  assign n28287 = ~n21589 ;
  assign n21590 = x[5] & n28287 ;
  assign n21591 = n27813 & n21589 ;
  assign n21592 = n21590 | n21591 ;
  assign n19257 = n19254 & n19256 ;
  assign n20334 = n19254 | n19256 ;
  assign n28288 = ~n19257 ;
  assign n20335 = n28288 & n20334 ;
  assign n28289 = ~n19440 ;
  assign n20336 = n28289 & n20335 ;
  assign n28290 = ~n20335 ;
  assign n20566 = n19440 & n28290 ;
  assign n20567 = n20336 | n20566 ;
  assign n20568 = n20565 & n20567 ;
  assign n21202 = n20568 | n21201 ;
  assign n12701 = n1741 & n12695 ;
  assign n12654 = x[77] & n12633 ;
  assign n14358 = x[78] & n13533 ;
  assign n19235 = n12654 | n14358 ;
  assign n19236 = x[79] & n12631 ;
  assign n19237 = n19235 | n19236 ;
  assign n19238 = n12701 | n19237 ;
  assign n28291 = ~n19238 ;
  assign n19239 = x[11] & n28291 ;
  assign n19240 = n27892 & n19238 ;
  assign n19241 = n19239 | n19240 ;
  assign n28292 = ~n17075 ;
  assign n17776 = n28292 & n17774 ;
  assign n28293 = ~n17774 ;
  assign n18011 = n17075 & n28293 ;
  assign n18012 = n17776 | n18011 ;
  assign n18013 = n18010 & n18012 ;
  assign n18155 = n18013 | n18154 ;
  assign n10559 = n2750 & n10542 ;
  assign n10529 = x[74] & n10481 ;
  assign n11880 = x[75] & n11232 ;
  assign n17994 = n10529 | n11880 ;
  assign n17995 = x[76] & n10479 ;
  assign n17996 = n17994 | n17995 ;
  assign n17997 = n10559 | n17996 ;
  assign n28294 = ~n17997 ;
  assign n17998 = x[14] & n28294 ;
  assign n17999 = n27956 & n17997 ;
  assign n18000 = n17998 | n17999 ;
  assign n7182 = n5976 & n7162 ;
  assign n7101 = x[68] & n7100 ;
  assign n7673 = x[69] & n7647 ;
  assign n16043 = n7101 | n7673 ;
  assign n16044 = x[70] & n7098 ;
  assign n16045 = n16043 | n16044 ;
  assign n16046 = n7182 | n16045 ;
  assign n28295 = ~n16046 ;
  assign n16047 = x[20] & n28295 ;
  assign n16048 = n28114 & n16046 ;
  assign n16049 = n16047 | n16048 ;
  assign n27330 = x[23] & x[24] ;
  assign n318 = x[23] | x[24] ;
  assign n28296 = ~n27330 ;
  assign n319 = n28296 & n318 ;
  assign n14076 = x[64] & n319 ;
  assign n15025 = n14076 & n28259 ;
  assign n28297 = ~n14076 ;
  assign n15026 = n28297 & n15024 ;
  assign n15027 = n15025 | n15026 ;
  assign n6508 = n5302 & n6494 ;
  assign n5245 = x[65] & n5240 ;
  assign n6222 = x[66] & n6179 ;
  assign n15028 = n5245 | n6222 ;
  assign n15029 = x[67] & n5238 ;
  assign n15030 = n15028 | n15029 ;
  assign n15031 = n6508 | n15030 ;
  assign n28298 = ~n15031 ;
  assign n15032 = x[23] & n28298 ;
  assign n15033 = n28221 & n15031 ;
  assign n15034 = n15032 | n15033 ;
  assign n28299 = ~n15034 ;
  assign n15035 = n15027 & n28299 ;
  assign n28300 = ~n15027 ;
  assign n16050 = n28300 & n15034 ;
  assign n16051 = n15035 | n16050 ;
  assign n28301 = ~n16049 ;
  assign n16052 = n28301 & n16051 ;
  assign n28302 = ~n16051 ;
  assign n16115 = n16049 & n28302 ;
  assign n16116 = n16052 | n16115 ;
  assign n16117 = n16114 & n16116 ;
  assign n16962 = n16114 | n16116 ;
  assign n28303 = ~n16117 ;
  assign n16963 = n28303 & n16962 ;
  assign n8710 = n3733 & n8706 ;
  assign n8668 = x[71] & n8645 ;
  assign n9898 = x[72] & n9278 ;
  assign n16964 = n8668 | n9898 ;
  assign n16965 = x[73] & n8643 ;
  assign n16966 = n16964 | n16965 ;
  assign n16967 = n8710 | n16966 ;
  assign n28304 = ~n16967 ;
  assign n16968 = x[17] & n28304 ;
  assign n16969 = n28039 & n16967 ;
  assign n16970 = n16968 | n16969 ;
  assign n16971 = n16963 & n16970 ;
  assign n17079 = n16963 | n16970 ;
  assign n28305 = ~n16971 ;
  assign n17080 = n28305 & n17079 ;
  assign n16984 = n16975 & n16982 ;
  assign n17777 = n16984 | n17775 ;
  assign n28306 = ~n17777 ;
  assign n17778 = n17080 & n28306 ;
  assign n28307 = ~n17080 ;
  assign n18001 = n28307 & n17777 ;
  assign n18002 = n17778 | n18001 ;
  assign n18003 = n18000 & n18002 ;
  assign n18156 = n18000 | n18002 ;
  assign n28308 = ~n18003 ;
  assign n19103 = n28308 & n18156 ;
  assign n28309 = ~n18155 ;
  assign n19105 = n28309 & n19103 ;
  assign n28310 = ~n19103 ;
  assign n19242 = n18155 & n28310 ;
  assign n19243 = n19105 | n19242 ;
  assign n19244 = n19241 & n19243 ;
  assign n19246 = n19241 | n19243 ;
  assign n28311 = ~n19244 ;
  assign n19247 = n28311 & n19246 ;
  assign n20373 = n19437 & n20371 ;
  assign n20374 = n19436 | n20373 ;
  assign n20375 = n20335 & n20374 ;
  assign n20376 = n19257 | n20375 ;
  assign n28312 = ~n20376 ;
  assign n20377 = n19247 & n28312 ;
  assign n28313 = ~n19247 ;
  assign n20549 = n28313 & n20376 ;
  assign n20550 = n20377 | n20549 ;
  assign n15319 = n1003 & n15308 ;
  assign n15255 = x[80] & n15246 ;
  assign n17321 = x[81] & n16288 ;
  assign n20551 = n15255 | n17321 ;
  assign n20552 = x[82] & n15244 ;
  assign n20553 = n20551 | n20552 ;
  assign n20554 = n15319 | n20553 ;
  assign n28314 = ~n20554 ;
  assign n20555 = x[8] & n28314 ;
  assign n20556 = n27845 & n20554 ;
  assign n20557 = n20555 | n20556 ;
  assign n20558 = n20550 & n20557 ;
  assign n28315 = ~n19241 ;
  assign n19245 = n28315 & n19243 ;
  assign n28316 = ~n19243 ;
  assign n20332 = n19241 & n28316 ;
  assign n20333 = n19245 | n20332 ;
  assign n20378 = n20333 | n20376 ;
  assign n20379 = n20333 & n20376 ;
  assign n28317 = ~n20379 ;
  assign n20800 = n20378 & n28317 ;
  assign n20801 = n20557 | n20800 ;
  assign n28318 = ~n20558 ;
  assign n21203 = n28318 & n20801 ;
  assign n21204 = n21202 & n21203 ;
  assign n21593 = n21202 | n21203 ;
  assign n28319 = ~n21204 ;
  assign n21594 = n28319 & n21593 ;
  assign n28320 = ~n21592 ;
  assign n21892 = n28320 & n21594 ;
  assign n28321 = ~n21594 ;
  assign n22202 = n21592 & n28321 ;
  assign n22203 = n21892 | n22202 ;
  assign n28322 = ~n22203 ;
  assign n22204 = n21891 & n28322 ;
  assign n28323 = ~n21891 ;
  assign n22577 = n28323 & n22203 ;
  assign n22578 = n22204 | n22577 ;
  assign n525 = n523 & n524 ;
  assign n526 = n27636 | n525 ;
  assign n26308 = x[87] & x[88] ;
  assign n527 = x[87] | x[88] ;
  assign n28324 = ~n26308 ;
  assign n1717 = n28324 & n527 ;
  assign n1718 = n526 & n1717 ;
  assign n1719 = n526 | n1717 ;
  assign n28325 = ~n1718 ;
  assign n1720 = n28325 & n1719 ;
  assign n19673 = n1720 & n19656 ;
  assign n19737 = x[86] & n19723 ;
  assign n19849 = x[87] & n19829 ;
  assign n22579 = n19737 | n19849 ;
  assign n22580 = x[88] & n19655 ;
  assign n22581 = n22579 | n22580 ;
  assign n22582 = n19673 | n22581 ;
  assign n28326 = ~n22582 ;
  assign n22583 = x[2] & n28326 ;
  assign n22584 = n27790 & n22582 ;
  assign n22585 = n22583 | n22584 ;
  assign n28327 = ~n22585 ;
  assign n22586 = n22578 & n28327 ;
  assign n28328 = ~n22578 ;
  assign n22588 = n28328 & n22585 ;
  assign n22589 = n22586 | n22588 ;
  assign n22599 = n22590 & n22597 ;
  assign n22917 = n22599 | n22916 ;
  assign n22918 = n22589 & n22917 ;
  assign n27657 = n22589 | n22917 ;
  assign n28329 = ~n22918 ;
  assign n153 = n28329 & n27657 ;
  assign n22587 = n22578 & n22585 ;
  assign n22919 = n22587 | n22918 ;
  assign n528 = n526 & n527 ;
  assign n529 = n26308 | n528 ;
  assign n27634 = x[88] & x[89] ;
  assign n530 = x[88] | x[89] ;
  assign n28330 = ~n27634 ;
  assign n1450 = n28330 & n530 ;
  assign n28331 = ~n529 ;
  assign n1451 = n28331 & n1450 ;
  assign n28332 = ~n1450 ;
  assign n1452 = n529 & n28332 ;
  assign n1453 = n1451 | n1452 ;
  assign n19675 = n1453 & n19656 ;
  assign n19740 = x[87] & n19723 ;
  assign n19858 = x[88] & n19829 ;
  assign n22566 = n19740 | n19858 ;
  assign n22567 = x[89] & n19655 ;
  assign n22568 = n22566 | n22567 ;
  assign n22569 = n19675 | n22568 ;
  assign n28333 = ~n22569 ;
  assign n22570 = x[2] & n28333 ;
  assign n22571 = n27790 & n22569 ;
  assign n22572 = n22570 | n22571 ;
  assign n12702 = n1270 & n12695 ;
  assign n12637 = x[78] & n12633 ;
  assign n14360 = x[79] & n13533 ;
  assign n19220 = n12637 | n14360 ;
  assign n19221 = x[80] & n12631 ;
  assign n19222 = n19220 | n19221 ;
  assign n19223 = n12702 | n19222 ;
  assign n28334 = ~n19223 ;
  assign n19224 = x[11] & n28334 ;
  assign n19225 = n27892 & n19223 ;
  assign n19226 = n19224 | n19225 ;
  assign n16053 = n16049 & n16051 ;
  assign n16118 = n16053 | n16117 ;
  assign n7167 = n4790 & n7162 ;
  assign n7102 = x[69] & n7100 ;
  assign n7675 = x[70] & n7647 ;
  assign n16032 = n7102 | n7675 ;
  assign n16033 = x[71] & n7098 ;
  assign n16034 = n16032 | n16033 ;
  assign n16035 = n7167 | n16034 ;
  assign n28335 = ~n16035 ;
  assign n16036 = x[20] & n28335 ;
  assign n16037 = n28114 & n16035 ;
  assign n16038 = n16036 | n16037 ;
  assign n15036 = n15027 & n15034 ;
  assign n15037 = n14076 & n15024 ;
  assign n15038 = n15036 | n15037 ;
  assign n6422 = n5302 & n6408 ;
  assign n5300 = x[66] & n5240 ;
  assign n6228 = x[67] & n6179 ;
  assign n15039 = n5300 | n6228 ;
  assign n15040 = x[68] & n5238 ;
  assign n15041 = n15039 | n15040 ;
  assign n15042 = n6422 | n15041 ;
  assign n28336 = ~n15042 ;
  assign n15043 = x[23] & n28336 ;
  assign n15044 = n28221 & n15042 ;
  assign n15045 = n15043 | n15044 ;
  assign n14077 = x[26] & n28297 ;
  assign n27381 = x[25] & x[26] ;
  assign n320 = x[25] | x[26] ;
  assign n28337 = ~n27381 ;
  assign n321 = n28337 & n320 ;
  assign n452 = n319 & n321 ;
  assign n6438 = n452 & n6437 ;
  assign n28338 = ~n321 ;
  assign n322 = n319 & n28338 ;
  assign n14078 = x[65] & n322 ;
  assign n27429 = x[24] & x[25] ;
  assign n327 = x[24] | x[25] ;
  assign n28339 = ~n27429 ;
  assign n328 = n28339 & n327 ;
  assign n28340 = ~n319 ;
  assign n390 = n28340 & n328 ;
  assign n14079 = x[64] & n390 ;
  assign n14080 = n14078 | n14079 ;
  assign n14081 = n6438 | n14080 ;
  assign n28341 = ~n14081 ;
  assign n14082 = x[26] & n28341 ;
  assign n28342 = ~x[26] ;
  assign n14083 = n28342 & n14081 ;
  assign n14084 = n14082 | n14083 ;
  assign n28343 = ~n14084 ;
  assign n14085 = n14077 & n28343 ;
  assign n28344 = ~n14077 ;
  assign n15046 = n28344 & n14084 ;
  assign n15047 = n14085 | n15046 ;
  assign n28345 = ~n15045 ;
  assign n15048 = n28345 & n15047 ;
  assign n28346 = ~n15047 ;
  assign n15049 = n15045 & n28346 ;
  assign n15050 = n15048 | n15049 ;
  assign n28347 = ~n15050 ;
  assign n15051 = n15038 & n28347 ;
  assign n28348 = ~n15038 ;
  assign n16039 = n28348 & n15050 ;
  assign n16040 = n15051 | n16039 ;
  assign n16041 = n16038 | n16040 ;
  assign n16042 = n16038 & n16040 ;
  assign n28349 = ~n16042 ;
  assign n16119 = n16041 & n28349 ;
  assign n28350 = ~n16118 ;
  assign n16120 = n28350 & n16119 ;
  assign n28351 = ~n16119 ;
  assign n16948 = n16118 & n28351 ;
  assign n16949 = n16120 | n16948 ;
  assign n8733 = n2722 & n8706 ;
  assign n8693 = x[72] & n8645 ;
  assign n9870 = x[73] & n9278 ;
  assign n16950 = n8693 | n9870 ;
  assign n16951 = x[74] & n8643 ;
  assign n16952 = n16950 | n16951 ;
  assign n16953 = n8733 | n16952 ;
  assign n28352 = ~n16953 ;
  assign n16954 = x[17] & n28352 ;
  assign n16955 = n28039 & n16953 ;
  assign n16956 = n16954 | n16955 ;
  assign n28353 = ~n16956 ;
  assign n16959 = n16949 & n28353 ;
  assign n28354 = ~n16949 ;
  assign n16960 = n28354 & n16956 ;
  assign n16961 = n16959 | n16960 ;
  assign n17076 = n16975 | n16982 ;
  assign n17077 = n17075 & n17076 ;
  assign n17078 = n16984 | n17077 ;
  assign n17081 = n17078 & n17080 ;
  assign n17082 = n16971 | n17081 ;
  assign n17083 = n16961 | n17082 ;
  assign n17084 = n16961 & n17082 ;
  assign n28355 = ~n17084 ;
  assign n17979 = n17083 & n28355 ;
  assign n10570 = n1775 & n10542 ;
  assign n10489 = x[75] & n10481 ;
  assign n11924 = x[76] & n11232 ;
  assign n17980 = n10489 | n11924 ;
  assign n17981 = x[77] & n10479 ;
  assign n17982 = n17980 | n17981 ;
  assign n17983 = n10570 | n17982 ;
  assign n28356 = ~n17983 ;
  assign n17984 = x[14] & n28356 ;
  assign n17985 = n27956 & n17983 ;
  assign n17986 = n17984 | n17985 ;
  assign n28357 = ~n17986 ;
  assign n17987 = n17979 & n28357 ;
  assign n28358 = ~n17979 ;
  assign n19069 = n28358 & n17986 ;
  assign n19070 = n17987 | n19069 ;
  assign n19097 = n18142 & n19095 ;
  assign n19098 = n18037 | n19097 ;
  assign n19099 = n19071 & n19098 ;
  assign n19100 = n18024 | n19099 ;
  assign n19101 = n18152 & n19100 ;
  assign n19102 = n18013 | n19101 ;
  assign n19104 = n19102 & n19103 ;
  assign n19106 = n18003 | n19104 ;
  assign n19108 = n19070 | n19106 ;
  assign n19109 = n19070 & n19106 ;
  assign n28359 = ~n19109 ;
  assign n19230 = n19108 & n28359 ;
  assign n28360 = ~n19226 ;
  assign n19231 = n28360 & n19230 ;
  assign n28361 = ~n19230 ;
  assign n19233 = n19226 & n28361 ;
  assign n19234 = n19231 | n19233 ;
  assign n19443 = n19257 | n19442 ;
  assign n19444 = n19247 & n19443 ;
  assign n19445 = n19244 | n19444 ;
  assign n19446 = n19234 | n19445 ;
  assign n19447 = n19234 & n19445 ;
  assign n28362 = ~n19447 ;
  assign n20534 = n19446 & n28362 ;
  assign n15320 = n1057 & n15308 ;
  assign n15289 = x[81] & n15246 ;
  assign n17302 = x[82] & n16288 ;
  assign n20535 = n15289 | n17302 ;
  assign n20536 = x[83] & n15244 ;
  assign n20537 = n20535 | n20536 ;
  assign n20538 = n15320 | n20537 ;
  assign n28363 = ~n20538 ;
  assign n20539 = x[8] & n28363 ;
  assign n20540 = n27845 & n20538 ;
  assign n20541 = n20539 | n20540 ;
  assign n28364 = ~n20541 ;
  assign n20542 = n20534 & n28364 ;
  assign n28365 = ~n20534 ;
  assign n21140 = n28365 & n20541 ;
  assign n21141 = n20542 | n21140 ;
  assign n21142 = n20557 & n20800 ;
  assign n21205 = n21142 | n21204 ;
  assign n21206 = n21141 | n21205 ;
  assign n21208 = n21141 & n21205 ;
  assign n28366 = ~n21208 ;
  assign n21897 = n21206 & n28366 ;
  assign n18457 = n1213 & n18392 ;
  assign n18360 = x[84] & n18329 ;
  assign n18575 = x[85] & n18514 ;
  assign n21898 = n18360 | n18575 ;
  assign n21899 = x[86] & n18327 ;
  assign n21900 = n21898 | n21899 ;
  assign n21901 = n18457 | n21900 ;
  assign n28367 = ~n21901 ;
  assign n21902 = x[5] & n28367 ;
  assign n21903 = n27813 & n21901 ;
  assign n21904 = n21902 | n21903 ;
  assign n28368 = ~n21904 ;
  assign n21905 = n21897 & n28368 ;
  assign n28369 = ~n21897 ;
  assign n21906 = n28369 & n21904 ;
  assign n21907 = n21905 | n21906 ;
  assign n21595 = n21592 & n21594 ;
  assign n21604 = n21596 | n21603 ;
  assign n28370 = ~n21605 ;
  assign n22125 = n21604 & n28370 ;
  assign n28371 = ~n21617 ;
  assign n21618 = n21610 & n28371 ;
  assign n28372 = ~n21610 ;
  assign n22126 = n28372 & n21617 ;
  assign n22127 = n21618 | n22126 ;
  assign n22198 = n22127 & n22196 ;
  assign n22199 = n21619 | n22198 ;
  assign n22200 = n22125 & n22199 ;
  assign n22201 = n21605 | n22200 ;
  assign n22205 = n22201 & n22203 ;
  assign n22206 = n21595 | n22205 ;
  assign n28373 = ~n21907 ;
  assign n22207 = n28373 & n22206 ;
  assign n28374 = ~n22206 ;
  assign n22573 = n21907 & n28374 ;
  assign n22574 = n22207 | n22573 ;
  assign n28375 = ~n22572 ;
  assign n22575 = n28375 & n22574 ;
  assign n28376 = ~n22574 ;
  assign n22920 = n22572 & n28376 ;
  assign n22921 = n22575 | n22920 ;
  assign n22922 = n22919 | n22921 ;
  assign n22923 = n22919 & n22921 ;
  assign n28377 = ~n22923 ;
  assign n154 = n22922 & n28377 ;
  assign n22576 = n22572 & n22574 ;
  assign n22924 = n22576 | n22923 ;
  assign n19232 = n19226 & n19230 ;
  assign n20329 = n19226 | n19230 ;
  assign n28378 = ~n19232 ;
  assign n20330 = n28378 & n20329 ;
  assign n28379 = ~n19445 ;
  assign n20331 = n28379 & n20330 ;
  assign n28380 = ~n20330 ;
  assign n20544 = n19445 & n28380 ;
  assign n20545 = n20331 | n20544 ;
  assign n20546 = n20541 | n20545 ;
  assign n20547 = n20541 & n20545 ;
  assign n28381 = ~n20547 ;
  assign n20548 = n20546 & n28381 ;
  assign n28382 = ~n21205 ;
  assign n21207 = n20548 & n28382 ;
  assign n28383 = ~n20548 ;
  assign n21908 = n28383 & n21205 ;
  assign n21909 = n21207 | n21908 ;
  assign n21911 = n21904 & n21909 ;
  assign n21893 = n21592 | n21594 ;
  assign n28384 = ~n21595 ;
  assign n21894 = n28384 & n21893 ;
  assign n21895 = n21891 & n21894 ;
  assign n21896 = n21595 | n21895 ;
  assign n21912 = n21896 & n21907 ;
  assign n21913 = n21911 | n21912 ;
  assign n16957 = n16949 | n16956 ;
  assign n16958 = n16949 & n16956 ;
  assign n28385 = ~n16958 ;
  assign n17771 = n16957 & n28385 ;
  assign n28386 = ~n17082 ;
  assign n17772 = n28386 & n17771 ;
  assign n28387 = ~n17771 ;
  assign n17989 = n17082 & n28387 ;
  assign n17990 = n17772 | n17989 ;
  assign n17991 = n17986 | n17990 ;
  assign n17992 = n17986 & n17990 ;
  assign n28388 = ~n17992 ;
  assign n17993 = n17991 & n28388 ;
  assign n28389 = ~n19106 ;
  assign n19107 = n17993 & n28389 ;
  assign n28390 = ~n17993 ;
  assign n19227 = n28390 & n19106 ;
  assign n19228 = n19107 | n19227 ;
  assign n19229 = n19226 & n19228 ;
  assign n19448 = n19229 | n19447 ;
  assign n10549 = n2084 & n10542 ;
  assign n10490 = x[76] & n10481 ;
  assign n11923 = x[77] & n11232 ;
  assign n17969 = n10490 | n11923 ;
  assign n17970 = x[78] & n10479 ;
  assign n17971 = n17969 | n17970 ;
  assign n17972 = n10549 | n17971 ;
  assign n28391 = ~n17972 ;
  assign n17973 = x[14] & n28391 ;
  assign n17974 = n27956 & n17972 ;
  assign n17975 = n17973 | n17974 ;
  assign n17085 = n16958 | n17084 ;
  assign n8717 = n3289 & n8706 ;
  assign n8695 = x[73] & n8645 ;
  assign n9897 = x[74] & n9278 ;
  assign n16938 = n8695 | n9897 ;
  assign n16939 = x[75] & n8643 ;
  assign n16940 = n16938 | n16939 ;
  assign n16941 = n8717 | n16940 ;
  assign n28392 = ~n16941 ;
  assign n16942 = x[17] & n28392 ;
  assign n16943 = n28039 & n16941 ;
  assign n16944 = n16942 | n16943 ;
  assign n16121 = n16118 & n16119 ;
  assign n16122 = n16042 | n16121 ;
  assign n14086 = n14077 & n14084 ;
  assign n6474 = n452 & n6466 ;
  assign n329 = n28340 & n321 ;
  assign n28393 = ~n328 ;
  assign n330 = n28393 & n329 ;
  assign n331 = x[64] & n330 ;
  assign n447 = x[65] & n390 ;
  assign n14087 = n331 | n447 ;
  assign n14088 = x[66] & n322 ;
  assign n14089 = n14087 | n14088 ;
  assign n14090 = n6474 | n14089 ;
  assign n28394 = ~n14090 ;
  assign n14091 = x[26] & n28394 ;
  assign n14092 = n28342 & n14090 ;
  assign n14093 = n14091 | n14092 ;
  assign n14094 = n14086 | n14093 ;
  assign n14095 = n14086 & n14093 ;
  assign n28395 = ~n14095 ;
  assign n14996 = n14094 & n28395 ;
  assign n6393 = n5302 & n6379 ;
  assign n5286 = x[67] & n5240 ;
  assign n6280 = x[68] & n6179 ;
  assign n14997 = n5286 | n6280 ;
  assign n14998 = x[69] & n5238 ;
  assign n14999 = n14997 | n14998 ;
  assign n15000 = n6393 | n14999 ;
  assign n28396 = ~n15000 ;
  assign n15001 = x[23] & n28396 ;
  assign n15002 = n28221 & n15000 ;
  assign n15003 = n15001 | n15002 ;
  assign n15055 = n14996 | n15003 ;
  assign n15004 = n14996 & n15003 ;
  assign n15052 = n15038 & n15050 ;
  assign n15053 = n15045 & n15047 ;
  assign n15054 = n15052 | n15053 ;
  assign n15056 = n15054 & n15055 ;
  assign n15058 = n15004 | n15056 ;
  assign n28397 = ~n15058 ;
  assign n15059 = n15055 & n28397 ;
  assign n28398 = ~n15004 ;
  assign n15057 = n28398 & n15055 ;
  assign n28399 = ~n15057 ;
  assign n16021 = n15054 & n28399 ;
  assign n16022 = n15059 | n16021 ;
  assign n7184 = n3701 & n7162 ;
  assign n7103 = x[70] & n7100 ;
  assign n7681 = x[71] & n7647 ;
  assign n16023 = n7103 | n7681 ;
  assign n16024 = x[72] & n7098 ;
  assign n16025 = n16023 | n16024 ;
  assign n16026 = n7184 | n16025 ;
  assign n28400 = ~n16026 ;
  assign n16027 = x[20] & n28400 ;
  assign n16028 = n28114 & n16026 ;
  assign n16029 = n16027 | n16028 ;
  assign n16030 = n16022 | n16029 ;
  assign n16031 = n16022 & n16029 ;
  assign n28401 = ~n16031 ;
  assign n16425 = n16030 & n28401 ;
  assign n16426 = n16122 & n16425 ;
  assign n17086 = n16122 | n16425 ;
  assign n28402 = ~n16426 ;
  assign n17087 = n28402 & n17086 ;
  assign n17088 = n16944 & n17087 ;
  assign n17089 = n16944 | n17087 ;
  assign n28403 = ~n17088 ;
  assign n17090 = n28403 & n17089 ;
  assign n17091 = n17085 & n17090 ;
  assign n17976 = n17085 | n17090 ;
  assign n28404 = ~n17091 ;
  assign n17977 = n28404 & n17976 ;
  assign n28405 = ~n17975 ;
  assign n18161 = n28405 & n17977 ;
  assign n28406 = ~n17977 ;
  assign n18162 = n17975 & n28406 ;
  assign n18163 = n18161 | n18162 ;
  assign n19110 = n17992 | n19109 ;
  assign n28407 = ~n18163 ;
  assign n19111 = n28407 & n19110 ;
  assign n28408 = ~n19110 ;
  assign n19210 = n18163 & n28408 ;
  assign n19211 = n19111 | n19210 ;
  assign n12706 = n1029 & n12695 ;
  assign n12648 = x[79] & n12633 ;
  assign n14361 = x[80] & n13533 ;
  assign n19212 = n12648 | n14361 ;
  assign n19213 = x[81] & n12631 ;
  assign n19214 = n19212 | n19213 ;
  assign n19215 = n12706 | n19214 ;
  assign n28409 = ~n19215 ;
  assign n19216 = x[11] & n28409 ;
  assign n19217 = n27892 & n19215 ;
  assign n19218 = n19216 | n19217 ;
  assign n19219 = n19211 & n19218 ;
  assign n19449 = n19211 | n19218 ;
  assign n28410 = ~n19219 ;
  assign n19450 = n28410 & n19449 ;
  assign n19451 = n19448 & n19450 ;
  assign n20520 = n19448 | n19450 ;
  assign n28411 = ~n19451 ;
  assign n20521 = n28411 & n20520 ;
  assign n15321 = n1293 & n15308 ;
  assign n15278 = x[82] & n15246 ;
  assign n17283 = x[83] & n16288 ;
  assign n20522 = n15278 | n17283 ;
  assign n20523 = x[84] & n15244 ;
  assign n20524 = n20522 | n20523 ;
  assign n20525 = n15321 | n20524 ;
  assign n28412 = ~n20525 ;
  assign n20526 = x[8] & n28412 ;
  assign n20527 = n27845 & n20525 ;
  assign n20528 = n20526 | n20527 ;
  assign n28413 = ~n20528 ;
  assign n20531 = n20521 & n28413 ;
  assign n28414 = ~n20521 ;
  assign n20532 = n28414 & n20528 ;
  assign n20533 = n20531 | n20532 ;
  assign n20543 = n20534 & n20541 ;
  assign n20791 = n20789 & n20790 ;
  assign n20792 = n20578 | n20791 ;
  assign n20794 = n20565 & n20793 ;
  assign n20796 = n20565 | n20793 ;
  assign n28415 = ~n20794 ;
  assign n20797 = n28415 & n20796 ;
  assign n20798 = n20792 & n20797 ;
  assign n20799 = n20568 | n20798 ;
  assign n20802 = n20799 & n20801 ;
  assign n20803 = n20558 | n20802 ;
  assign n20804 = n20548 & n20803 ;
  assign n20805 = n20543 | n20804 ;
  assign n20806 = n20533 | n20805 ;
  assign n20807 = n20533 & n20805 ;
  assign n28416 = ~n20807 ;
  assign n21576 = n20806 & n28416 ;
  assign n18407 = n1522 & n18392 ;
  assign n18338 = x[85] & n18329 ;
  assign n18527 = x[86] & n18514 ;
  assign n21577 = n18338 | n18527 ;
  assign n21578 = x[87] & n18327 ;
  assign n21579 = n21577 | n21578 ;
  assign n21580 = n18407 | n21579 ;
  assign n28417 = ~n21580 ;
  assign n21581 = x[5] & n28417 ;
  assign n21582 = n27813 & n21580 ;
  assign n21583 = n21581 | n21582 ;
  assign n28418 = ~n21583 ;
  assign n21584 = n21576 & n28418 ;
  assign n28419 = ~n21576 ;
  assign n22212 = n28419 & n21583 ;
  assign n22213 = n21584 | n22212 ;
  assign n28420 = ~n22213 ;
  assign n22214 = n21913 & n28420 ;
  assign n28421 = ~n21913 ;
  assign n22555 = n28421 & n22213 ;
  assign n22556 = n22214 | n22555 ;
  assign n531 = n529 & n530 ;
  assign n532 = n27634 | n531 ;
  assign n26187 = x[89] & x[90] ;
  assign n533 = x[89] | x[90] ;
  assign n28422 = ~n26187 ;
  assign n1479 = n28422 & n533 ;
  assign n1480 = n532 & n1479 ;
  assign n1481 = n532 | n1479 ;
  assign n28423 = ~n1480 ;
  assign n1482 = n28423 & n1481 ;
  assign n19676 = n1482 & n19656 ;
  assign n19744 = x[88] & n19723 ;
  assign n19851 = x[89] & n19829 ;
  assign n22557 = n19744 | n19851 ;
  assign n22558 = x[90] & n19655 ;
  assign n22559 = n22557 | n22558 ;
  assign n22560 = n19676 | n22559 ;
  assign n28424 = ~n22560 ;
  assign n22561 = x[2] & n28424 ;
  assign n22562 = n27790 & n22560 ;
  assign n22563 = n22561 | n22562 ;
  assign n22564 = n22556 | n22563 ;
  assign n22565 = n22556 & n22563 ;
  assign n28425 = ~n22565 ;
  assign n22925 = n22564 & n28425 ;
  assign n22926 = n22924 & n22925 ;
  assign n27660 = n22924 | n22925 ;
  assign n28426 = ~n22926 ;
  assign n155 = n28426 & n27660 ;
  assign n22927 = n22565 | n22926 ;
  assign n21585 = n21576 & n21583 ;
  assign n20529 = n20521 | n20528 ;
  assign n20530 = n20521 & n20528 ;
  assign n28427 = ~n20530 ;
  assign n21138 = n20529 & n28427 ;
  assign n28428 = ~n20805 ;
  assign n21139 = n28428 & n21138 ;
  assign n28429 = ~n21138 ;
  assign n21914 = n20805 & n28429 ;
  assign n21915 = n21139 | n21914 ;
  assign n21916 = n21583 | n21915 ;
  assign n21917 = n21583 & n21915 ;
  assign n28430 = ~n21917 ;
  assign n21918 = n21916 & n28430 ;
  assign n21919 = n21913 & n21918 ;
  assign n21920 = n21585 | n21919 ;
  assign n18404 = n1720 & n18392 ;
  assign n18345 = x[86] & n18329 ;
  assign n18543 = x[87] & n18514 ;
  assign n21561 = n18345 | n18543 ;
  assign n21562 = x[88] & n18327 ;
  assign n21563 = n21561 | n21562 ;
  assign n21564 = n18404 | n21563 ;
  assign n28431 = ~n21564 ;
  assign n21565 = x[5] & n28431 ;
  assign n21566 = n27813 & n21564 ;
  assign n21567 = n21565 | n21566 ;
  assign n12707 = n1003 & n12695 ;
  assign n12640 = x[80] & n12633 ;
  assign n14364 = x[81] & n13533 ;
  assign n19197 = n12640 | n14364 ;
  assign n19198 = x[82] & n12631 ;
  assign n19199 = n19197 | n19198 ;
  assign n19200 = n12707 | n19199 ;
  assign n28432 = ~n19200 ;
  assign n19201 = x[11] & n28432 ;
  assign n19202 = n27892 & n19200 ;
  assign n19203 = n19201 | n19202 ;
  assign n10551 = n1741 & n10542 ;
  assign n10497 = x[77] & n10481 ;
  assign n11910 = x[78] & n11232 ;
  assign n17956 = n10497 | n11910 ;
  assign n17957 = x[79] & n10479 ;
  assign n17958 = n17956 | n17957 ;
  assign n17959 = n10551 | n17958 ;
  assign n28433 = ~n17959 ;
  assign n17960 = x[14] & n28433 ;
  assign n17961 = n27956 & n17959 ;
  assign n17962 = n17960 | n17961 ;
  assign n28434 = ~n16122 ;
  assign n16427 = n28434 & n16425 ;
  assign n28435 = ~n16425 ;
  assign n16945 = n16122 & n28435 ;
  assign n16946 = n16427 | n16945 ;
  assign n16947 = n16944 & n16946 ;
  assign n17092 = n16947 | n17091 ;
  assign n8734 = n2750 & n8706 ;
  assign n8649 = x[74] & n8645 ;
  assign n9896 = x[75] & n9278 ;
  assign n16928 = n8649 | n9896 ;
  assign n16929 = x[76] & n8643 ;
  assign n16930 = n16928 | n16929 ;
  assign n16931 = n8734 | n16930 ;
  assign n28436 = ~n16931 ;
  assign n16932 = x[17] & n28436 ;
  assign n16933 = n28039 & n16931 ;
  assign n16934 = n16932 | n16933 ;
  assign n7163 = n3733 & n7162 ;
  assign n7152 = x[71] & n7100 ;
  assign n7677 = x[72] & n7647 ;
  assign n16013 = n7152 | n7677 ;
  assign n16014 = x[73] & n7098 ;
  assign n16015 = n16013 | n16014 ;
  assign n16016 = n7163 | n16015 ;
  assign n28437 = ~n16016 ;
  assign n16017 = x[20] & n28437 ;
  assign n16018 = n28114 & n16016 ;
  assign n16019 = n16017 | n16018 ;
  assign n5978 = n5302 & n5976 ;
  assign n5241 = x[68] & n5240 ;
  assign n6236 = x[69] & n6179 ;
  assign n14985 = n5241 | n6236 ;
  assign n14986 = x[70] & n5238 ;
  assign n14987 = n14985 | n14986 ;
  assign n14988 = n5978 | n14987 ;
  assign n28438 = ~n14988 ;
  assign n14989 = x[23] & n28438 ;
  assign n14990 = n28221 & n14988 ;
  assign n14991 = n14989 | n14990 ;
  assign n27760 = x[26] & x[27] ;
  assign n4500 = x[26] | x[27] ;
  assign n28439 = ~n27760 ;
  assign n4501 = n28439 & n4500 ;
  assign n13298 = x[64] & n4501 ;
  assign n14096 = n13298 & n28395 ;
  assign n28440 = ~n13298 ;
  assign n14097 = n28440 & n14095 ;
  assign n14098 = n14096 | n14097 ;
  assign n6495 = n452 & n6494 ;
  assign n332 = x[65] & n330 ;
  assign n437 = x[66] & n390 ;
  assign n14099 = n332 | n437 ;
  assign n14100 = x[67] & n322 ;
  assign n14101 = n14099 | n14100 ;
  assign n14102 = n6495 | n14101 ;
  assign n28441 = ~n14102 ;
  assign n14103 = x[26] & n28441 ;
  assign n14104 = n28342 & n14102 ;
  assign n14105 = n14103 | n14104 ;
  assign n28442 = ~n14105 ;
  assign n14106 = n14098 & n28442 ;
  assign n28443 = ~n14098 ;
  assign n14992 = n28443 & n14105 ;
  assign n14993 = n14106 | n14992 ;
  assign n28444 = ~n14991 ;
  assign n14994 = n28444 & n14993 ;
  assign n28445 = ~n14993 ;
  assign n15060 = n14991 & n28445 ;
  assign n15061 = n14994 | n15060 ;
  assign n28446 = ~n15061 ;
  assign n15748 = n15058 & n28446 ;
  assign n16125 = n28397 & n15061 ;
  assign n16126 = n15748 | n16125 ;
  assign n16127 = n16019 & n16126 ;
  assign n15062 = n15058 | n15061 ;
  assign n15063 = n15058 & n15061 ;
  assign n28447 = ~n15063 ;
  assign n16012 = n15062 & n28447 ;
  assign n16128 = n16012 | n16019 ;
  assign n28448 = ~n16127 ;
  assign n16129 = n28448 & n16128 ;
  assign n16428 = n16031 | n16426 ;
  assign n28449 = ~n16428 ;
  assign n16429 = n16129 & n28449 ;
  assign n28450 = ~n16129 ;
  assign n16935 = n28450 & n16428 ;
  assign n16936 = n16429 | n16935 ;
  assign n16937 = n16934 & n16936 ;
  assign n17093 = n16934 | n16936 ;
  assign n28451 = ~n16937 ;
  assign n17785 = n28451 & n17093 ;
  assign n28452 = ~n17092 ;
  assign n17787 = n28452 & n17785 ;
  assign n28453 = ~n17785 ;
  assign n17963 = n17092 & n28453 ;
  assign n17964 = n17787 | n17963 ;
  assign n28454 = ~n17962 ;
  assign n17966 = n28454 & n17964 ;
  assign n28455 = ~n17964 ;
  assign n19067 = n17962 & n28455 ;
  assign n19068 = n17966 | n19067 ;
  assign n17978 = n17975 & n17977 ;
  assign n19112 = n17975 | n17977 ;
  assign n28456 = ~n17978 ;
  assign n19113 = n28456 & n19112 ;
  assign n19114 = n19110 & n19113 ;
  assign n19115 = n17978 | n19114 ;
  assign n19117 = n19068 | n19115 ;
  assign n19118 = n19068 & n19115 ;
  assign n28457 = ~n19118 ;
  assign n19206 = n19117 & n28457 ;
  assign n28458 = ~n19203 ;
  assign n19207 = n28458 & n19206 ;
  assign n28459 = ~n19206 ;
  assign n19208 = n19203 & n28459 ;
  assign n19209 = n19207 | n19208 ;
  assign n19452 = n19219 | n19451 ;
  assign n19453 = n19209 | n19452 ;
  assign n19454 = n19209 & n19452 ;
  assign n28460 = ~n19454 ;
  assign n20505 = n19453 & n28460 ;
  assign n15323 = n1239 & n15308 ;
  assign n15270 = x[83] & n15246 ;
  assign n17332 = x[84] & n16288 ;
  assign n20506 = n15270 | n17332 ;
  assign n20507 = x[85] & n15244 ;
  assign n20508 = n20506 | n20507 ;
  assign n20509 = n15323 | n20508 ;
  assign n28461 = ~n20509 ;
  assign n20510 = x[8] & n28461 ;
  assign n20511 = n27845 & n20509 ;
  assign n20512 = n20510 | n20511 ;
  assign n28462 = ~n20512 ;
  assign n20513 = n20505 & n28462 ;
  assign n28463 = ~n20505 ;
  assign n21136 = n28463 & n20512 ;
  assign n21137 = n20513 | n21136 ;
  assign n21209 = n20547 | n21208 ;
  assign n21210 = n21138 & n21209 ;
  assign n21211 = n20530 | n21210 ;
  assign n21213 = n21137 | n21211 ;
  assign n21214 = n21137 & n21211 ;
  assign n28464 = ~n21214 ;
  assign n21571 = n21213 & n28464 ;
  assign n21573 = n21567 & n21571 ;
  assign n22122 = n21567 | n21571 ;
  assign n28465 = ~n21573 ;
  assign n22123 = n28465 & n22122 ;
  assign n28466 = ~n21920 ;
  assign n22124 = n28466 & n22123 ;
  assign n28467 = ~n22123 ;
  assign n22544 = n21920 & n28467 ;
  assign n22545 = n22124 | n22544 ;
  assign n534 = n532 & n533 ;
  assign n535 = n26187 | n534 ;
  assign n27633 = x[90] & x[91] ;
  assign n536 = x[90] | x[91] ;
  assign n28468 = ~n27633 ;
  assign n2043 = n28468 & n536 ;
  assign n2044 = n535 | n2043 ;
  assign n2045 = n535 & n2043 ;
  assign n28469 = ~n2045 ;
  assign n2046 = n2044 & n28469 ;
  assign n19708 = n2046 & n19656 ;
  assign n19753 = x[89] & n19723 ;
  assign n19854 = x[90] & n19829 ;
  assign n22546 = n19753 | n19854 ;
  assign n22547 = x[91] & n19655 ;
  assign n22548 = n22546 | n22547 ;
  assign n22549 = n19708 | n22548 ;
  assign n28470 = ~n22549 ;
  assign n22550 = x[2] & n28470 ;
  assign n22551 = n27790 & n22549 ;
  assign n22552 = n22550 | n22551 ;
  assign n22553 = n22545 | n22552 ;
  assign n22554 = n22545 & n22552 ;
  assign n28471 = ~n22554 ;
  assign n22928 = n22553 & n28471 ;
  assign n22929 = n22927 | n22928 ;
  assign n22930 = n22927 & n22928 ;
  assign n28472 = ~n22930 ;
  assign n156 = n22929 & n28472 ;
  assign n22931 = n22554 | n22930 ;
  assign n18405 = n1453 & n18392 ;
  assign n18339 = x[87] & n18329 ;
  assign n18525 = x[88] & n18514 ;
  assign n21546 = n18339 | n18525 ;
  assign n21547 = x[89] & n18327 ;
  assign n21548 = n21546 | n21547 ;
  assign n21549 = n18405 | n21548 ;
  assign n28473 = ~n21549 ;
  assign n21550 = x[5] & n28473 ;
  assign n21551 = n27813 & n21549 ;
  assign n21552 = n21550 | n21551 ;
  assign n15333 = n1213 & n15308 ;
  assign n15303 = x[84] & n15246 ;
  assign n17286 = x[85] & n16288 ;
  assign n20492 = n15303 | n17286 ;
  assign n20493 = x[86] & n15244 ;
  assign n20494 = n20492 | n20493 ;
  assign n20495 = n15333 | n20494 ;
  assign n28474 = ~n20495 ;
  assign n20496 = x[8] & n28474 ;
  assign n20497 = n27845 & n20495 ;
  assign n20498 = n20496 | n20497 ;
  assign n10552 = n1270 & n10542 ;
  assign n10491 = x[78] & n10481 ;
  assign n11879 = x[79] & n11232 ;
  assign n17943 = n10491 | n11879 ;
  assign n17944 = x[80] & n10479 ;
  assign n17945 = n17943 | n17944 ;
  assign n17946 = n10552 | n17945 ;
  assign n28475 = ~n17946 ;
  assign n17947 = x[14] & n28475 ;
  assign n17948 = n27956 & n17946 ;
  assign n17949 = n17947 | n17948 ;
  assign n14995 = n14991 & n14993 ;
  assign n15064 = n14995 | n15063 ;
  assign n5331 = n4790 & n5302 ;
  assign n5257 = x[69] & n5240 ;
  assign n6248 = x[70] & n6179 ;
  assign n14975 = n5257 | n6248 ;
  assign n14976 = x[71] & n5238 ;
  assign n14977 = n14975 | n14976 ;
  assign n14978 = n5331 | n14977 ;
  assign n28476 = ~n14978 ;
  assign n14979 = x[23] & n28476 ;
  assign n14980 = n28221 & n14978 ;
  assign n14981 = n14979 | n14980 ;
  assign n14107 = n14098 & n14105 ;
  assign n14108 = n13298 & n14095 ;
  assign n14109 = n14107 | n14108 ;
  assign n6409 = n452 & n6408 ;
  assign n370 = x[66] & n330 ;
  assign n448 = x[67] & n390 ;
  assign n14110 = n370 | n448 ;
  assign n14111 = x[68] & n322 ;
  assign n14112 = n14110 | n14111 ;
  assign n14113 = n6409 | n14112 ;
  assign n28477 = ~n14113 ;
  assign n14114 = x[26] & n28477 ;
  assign n14115 = n28342 & n14113 ;
  assign n14116 = n14114 | n14115 ;
  assign n13299 = x[29] & n28440 ;
  assign n27761 = x[28] & x[29] ;
  assign n4502 = x[28] | x[29] ;
  assign n28478 = ~n27761 ;
  assign n4503 = n28478 & n4502 ;
  assign n4632 = n4501 & n4503 ;
  assign n6445 = n4632 & n6437 ;
  assign n28479 = ~n4503 ;
  assign n4504 = n4501 & n28479 ;
  assign n13300 = x[65] & n4504 ;
  assign n27763 = x[27] & x[28] ;
  assign n4511 = x[27] | x[28] ;
  assign n28480 = ~n27763 ;
  assign n4512 = n28480 & n4511 ;
  assign n28481 = ~n4501 ;
  assign n4572 = n28481 & n4512 ;
  assign n13301 = x[64] & n4572 ;
  assign n13302 = n13300 | n13301 ;
  assign n13303 = n6445 | n13302 ;
  assign n28482 = ~n13303 ;
  assign n13304 = x[29] & n28482 ;
  assign n28483 = ~x[29] ;
  assign n13305 = n28483 & n13303 ;
  assign n13306 = n13304 | n13305 ;
  assign n28484 = ~n13306 ;
  assign n13307 = n13299 & n28484 ;
  assign n28485 = ~n13299 ;
  assign n14117 = n28485 & n13306 ;
  assign n14118 = n13307 | n14117 ;
  assign n28486 = ~n14116 ;
  assign n14119 = n28486 & n14118 ;
  assign n28487 = ~n14118 ;
  assign n14120 = n14116 & n28487 ;
  assign n14121 = n14119 | n14120 ;
  assign n28488 = ~n14121 ;
  assign n14122 = n14109 & n28488 ;
  assign n28489 = ~n14109 ;
  assign n14982 = n28489 & n14121 ;
  assign n14983 = n14122 | n14982 ;
  assign n14984 = n14981 & n14983 ;
  assign n15065 = n14981 | n14983 ;
  assign n28490 = ~n14984 ;
  assign n15066 = n28490 & n15065 ;
  assign n15067 = n15064 & n15066 ;
  assign n15998 = n15064 | n15066 ;
  assign n28491 = ~n15067 ;
  assign n15999 = n28491 & n15998 ;
  assign n7164 = n2722 & n7162 ;
  assign n7104 = x[72] & n7100 ;
  assign n7695 = x[73] & n7647 ;
  assign n16000 = n7104 | n7695 ;
  assign n16001 = x[74] & n7098 ;
  assign n16002 = n16000 | n16001 ;
  assign n16003 = n7164 | n16002 ;
  assign n28492 = ~n16003 ;
  assign n16004 = x[20] & n28492 ;
  assign n16005 = n28114 & n16003 ;
  assign n16006 = n16004 | n16005 ;
  assign n28493 = ~n16006 ;
  assign n16009 = n15999 & n28493 ;
  assign n28494 = ~n15999 ;
  assign n16010 = n28494 & n16006 ;
  assign n16011 = n16009 | n16010 ;
  assign n16020 = n16012 & n16019 ;
  assign n16123 = n16030 & n16122 ;
  assign n16124 = n16031 | n16123 ;
  assign n16130 = n16124 & n16129 ;
  assign n16131 = n16020 | n16130 ;
  assign n16132 = n16011 | n16131 ;
  assign n16133 = n16011 & n16131 ;
  assign n28495 = ~n16133 ;
  assign n16913 = n16132 & n28495 ;
  assign n8724 = n1775 & n8706 ;
  assign n8651 = x[75] & n8645 ;
  assign n9894 = x[76] & n9278 ;
  assign n16914 = n8651 | n9894 ;
  assign n16915 = x[77] & n8643 ;
  assign n16916 = n16914 | n16915 ;
  assign n16917 = n8724 | n16916 ;
  assign n28496 = ~n16917 ;
  assign n16918 = x[17] & n28496 ;
  assign n16919 = n28039 & n16917 ;
  assign n16920 = n16918 | n16919 ;
  assign n28497 = ~n16920 ;
  assign n16921 = n16913 & n28497 ;
  assign n28498 = ~n16913 ;
  assign n17769 = n28498 & n16920 ;
  assign n17770 = n16921 | n17769 ;
  assign n17779 = n17079 & n17777 ;
  assign n17780 = n16971 | n17779 ;
  assign n17781 = n17771 & n17780 ;
  assign n17782 = n16958 | n17781 ;
  assign n17783 = n17089 & n17782 ;
  assign n17784 = n16947 | n17783 ;
  assign n17786 = n17784 & n17785 ;
  assign n17788 = n16937 | n17786 ;
  assign n17790 = n17770 | n17788 ;
  assign n17791 = n17770 & n17788 ;
  assign n28499 = ~n17791 ;
  assign n17952 = n17790 & n28499 ;
  assign n28500 = ~n17949 ;
  assign n17953 = n28500 & n17952 ;
  assign n28501 = ~n17952 ;
  assign n17954 = n17949 & n28501 ;
  assign n17955 = n17953 | n17954 ;
  assign n17965 = n17962 & n17964 ;
  assign n17967 = n17962 | n17964 ;
  assign n28502 = ~n17965 ;
  assign n17968 = n28502 & n17967 ;
  assign n17988 = n17979 & n17986 ;
  assign n18157 = n18155 & n18156 ;
  assign n18158 = n18003 | n18157 ;
  assign n18159 = n17993 & n18158 ;
  assign n18160 = n17988 | n18159 ;
  assign n18164 = n18160 & n18163 ;
  assign n18165 = n17978 | n18164 ;
  assign n18166 = n17968 & n18165 ;
  assign n18167 = n17965 | n18166 ;
  assign n18168 = n17955 | n18167 ;
  assign n18169 = n17955 & n18167 ;
  assign n28503 = ~n18169 ;
  assign n19180 = n18168 & n28503 ;
  assign n12718 = n1057 & n12695 ;
  assign n12641 = x[81] & n12633 ;
  assign n14395 = x[82] & n13533 ;
  assign n19181 = n12641 | n14395 ;
  assign n19182 = x[83] & n12631 ;
  assign n19183 = n19181 | n19182 ;
  assign n19184 = n12718 | n19183 ;
  assign n28504 = ~n19184 ;
  assign n19185 = x[11] & n28504 ;
  assign n19186 = n27892 & n19184 ;
  assign n19187 = n19185 | n19186 ;
  assign n28505 = ~n19187 ;
  assign n19188 = n19180 & n28505 ;
  assign n28506 = ~n19180 ;
  assign n20324 = n28506 & n19187 ;
  assign n20325 = n19188 | n20324 ;
  assign n20326 = n19203 & n19206 ;
  assign n28507 = ~n19115 ;
  assign n19116 = n17968 & n28507 ;
  assign n28508 = ~n17968 ;
  assign n19195 = n28508 & n19115 ;
  assign n19196 = n19116 | n19195 ;
  assign n19204 = n19196 | n19203 ;
  assign n19205 = n19196 & n19203 ;
  assign n28509 = ~n19205 ;
  assign n20327 = n19204 & n28509 ;
  assign n20380 = n19244 | n20379 ;
  assign n20381 = n20330 & n20380 ;
  assign n20382 = n19229 | n20381 ;
  assign n20383 = n19449 & n20382 ;
  assign n20384 = n19219 | n20383 ;
  assign n20385 = n20327 & n20384 ;
  assign n20386 = n20326 | n20385 ;
  assign n20388 = n20325 | n20386 ;
  assign n20389 = n20325 & n20386 ;
  assign n28510 = ~n20389 ;
  assign n20501 = n20388 & n28510 ;
  assign n28511 = ~n20498 ;
  assign n20502 = n28511 & n20501 ;
  assign n28512 = ~n20501 ;
  assign n20503 = n20498 & n28512 ;
  assign n20504 = n20502 | n20503 ;
  assign n20514 = n20505 & n20512 ;
  assign n28513 = ~n19452 ;
  assign n20328 = n28513 & n20327 ;
  assign n28514 = ~n20327 ;
  assign n20515 = n19452 & n28514 ;
  assign n20516 = n20328 | n20515 ;
  assign n20517 = n20512 | n20516 ;
  assign n20518 = n20512 & n20516 ;
  assign n28515 = ~n20518 ;
  assign n20519 = n20517 & n28515 ;
  assign n20808 = n20530 | n20807 ;
  assign n20809 = n20519 & n20808 ;
  assign n20810 = n20514 | n20809 ;
  assign n20811 = n20504 | n20810 ;
  assign n20812 = n20504 & n20810 ;
  assign n28516 = ~n20812 ;
  assign n21556 = n20811 & n28516 ;
  assign n21557 = n21552 & n21556 ;
  assign n21559 = n21552 | n21556 ;
  assign n28517 = ~n21557 ;
  assign n21560 = n28517 & n21559 ;
  assign n28518 = ~n21211 ;
  assign n21212 = n20519 & n28518 ;
  assign n28519 = ~n20519 ;
  assign n21568 = n28519 & n21211 ;
  assign n21569 = n21212 | n21568 ;
  assign n21570 = n21567 & n21569 ;
  assign n21910 = n21904 | n21909 ;
  assign n28520 = ~n21911 ;
  assign n22208 = n21910 & n28520 ;
  assign n22209 = n22206 & n22208 ;
  assign n22210 = n21897 & n21904 ;
  assign n22211 = n22209 | n22210 ;
  assign n22215 = n22211 & n22213 ;
  assign n22216 = n21917 | n22215 ;
  assign n22217 = n22123 & n22216 ;
  assign n22218 = n21570 | n22217 ;
  assign n28521 = ~n22218 ;
  assign n22219 = n21560 & n28521 ;
  assign n28522 = ~n21560 ;
  assign n22533 = n28522 & n22218 ;
  assign n22534 = n22219 | n22533 ;
  assign n537 = n535 & n536 ;
  assign n538 = n27633 | n537 ;
  assign n26068 = x[91] & x[92] ;
  assign n539 = x[91] | x[92] ;
  assign n28523 = ~n26068 ;
  assign n1838 = n28523 & n539 ;
  assign n1839 = n538 & n1838 ;
  assign n1840 = n538 | n1838 ;
  assign n28524 = ~n1839 ;
  assign n1841 = n28524 & n1840 ;
  assign n19666 = n1841 & n19656 ;
  assign n19745 = x[90] & n19723 ;
  assign n19860 = x[91] & n19829 ;
  assign n22535 = n19745 | n19860 ;
  assign n22536 = x[92] & n19655 ;
  assign n22537 = n22535 | n22536 ;
  assign n22538 = n19666 | n22537 ;
  assign n28525 = ~n22538 ;
  assign n22539 = x[2] & n28525 ;
  assign n22540 = n27790 & n22538 ;
  assign n22541 = n22539 | n22540 ;
  assign n22542 = n22534 | n22541 ;
  assign n22543 = n22534 & n22541 ;
  assign n28526 = ~n22543 ;
  assign n22932 = n22542 & n28526 ;
  assign n22933 = n22931 & n22932 ;
  assign n27663 = n22931 | n22932 ;
  assign n28527 = ~n22933 ;
  assign n157 = n28527 & n27663 ;
  assign n18430 = n1482 & n18392 ;
  assign n18341 = x[88] & n18329 ;
  assign n18528 = x[89] & n18514 ;
  assign n21536 = n18341 | n18528 ;
  assign n21537 = x[90] & n18327 ;
  assign n21538 = n21536 | n21537 ;
  assign n21539 = n18430 | n21538 ;
  assign n28528 = ~n21539 ;
  assign n21540 = x[5] & n28528 ;
  assign n21541 = n27813 & n21539 ;
  assign n21542 = n21540 | n21541 ;
  assign n16007 = n15999 | n16006 ;
  assign n16008 = n15999 & n16006 ;
  assign n28529 = ~n16008 ;
  assign n16423 = n16007 & n28529 ;
  assign n28530 = ~n16131 ;
  assign n16424 = n28530 & n16423 ;
  assign n28531 = ~n16423 ;
  assign n16923 = n16131 & n28531 ;
  assign n16924 = n16424 | n16923 ;
  assign n16925 = n16920 | n16924 ;
  assign n16926 = n16920 & n16924 ;
  assign n28532 = ~n16926 ;
  assign n16927 = n16925 & n28532 ;
  assign n28533 = ~n17788 ;
  assign n17789 = n16927 & n28533 ;
  assign n28534 = ~n16927 ;
  assign n17941 = n28534 & n17788 ;
  assign n17942 = n17789 | n17941 ;
  assign n17950 = n17942 | n17949 ;
  assign n17951 = n17942 & n17949 ;
  assign n28535 = ~n17951 ;
  assign n19065 = n17950 & n28535 ;
  assign n28536 = ~n18167 ;
  assign n19066 = n28536 & n19065 ;
  assign n28537 = ~n19065 ;
  assign n19190 = n18167 & n28537 ;
  assign n19191 = n19066 | n19190 ;
  assign n19193 = n19187 & n19191 ;
  assign n20390 = n19193 | n20389 ;
  assign n10553 = n1029 & n10542 ;
  assign n10525 = x[79] & n10481 ;
  assign n11918 = x[80] & n11232 ;
  assign n17927 = n10525 | n11918 ;
  assign n17928 = x[81] & n10479 ;
  assign n17929 = n17927 | n17928 ;
  assign n17930 = n10553 | n17929 ;
  assign n28538 = ~n17930 ;
  assign n17931 = x[14] & n28538 ;
  assign n17932 = n27956 & n17930 ;
  assign n17933 = n17931 | n17932 ;
  assign n16922 = n16913 & n16920 ;
  assign n17094 = n17092 & n17093 ;
  assign n17095 = n16937 | n17094 ;
  assign n17096 = n16927 & n17095 ;
  assign n17097 = n16922 | n17096 ;
  assign n8714 = n2084 & n8706 ;
  assign n8653 = x[76] & n8645 ;
  assign n9860 = x[77] & n9278 ;
  assign n16900 = n8653 | n9860 ;
  assign n16901 = x[78] & n8643 ;
  assign n16902 = n16900 | n16901 ;
  assign n16903 = n8714 | n16902 ;
  assign n28539 = ~n16903 ;
  assign n16904 = x[17] & n28539 ;
  assign n16905 = n28039 & n16903 ;
  assign n16906 = n16904 | n16905 ;
  assign n16134 = n16008 | n16133 ;
  assign n7165 = n3289 & n7162 ;
  assign n7105 = x[73] & n7100 ;
  assign n7678 = x[74] & n7647 ;
  assign n15988 = n7105 | n7678 ;
  assign n15989 = x[75] & n7098 ;
  assign n15990 = n15988 | n15989 ;
  assign n15991 = n7165 | n15990 ;
  assign n28540 = ~n15991 ;
  assign n15992 = x[20] & n28540 ;
  assign n15993 = n28114 & n15991 ;
  assign n15994 = n15992 | n15993 ;
  assign n15068 = n14984 | n15067 ;
  assign n13308 = n13299 & n13306 ;
  assign n6478 = n4632 & n6466 ;
  assign n4513 = n28481 & n4503 ;
  assign n28541 = ~n4512 ;
  assign n4514 = n28541 & n4513 ;
  assign n4560 = x[64] & n4514 ;
  assign n4611 = x[65] & n4572 ;
  assign n13309 = n4560 | n4611 ;
  assign n13310 = x[66] & n4504 ;
  assign n13311 = n13309 | n13310 ;
  assign n13312 = n6478 | n13311 ;
  assign n28542 = ~n13312 ;
  assign n13313 = x[29] & n28542 ;
  assign n13314 = n28483 & n13312 ;
  assign n13315 = n13313 | n13314 ;
  assign n13316 = n13308 | n13315 ;
  assign n13317 = n13308 & n13315 ;
  assign n28543 = ~n13317 ;
  assign n14067 = n13316 & n28543 ;
  assign n6382 = n452 & n6379 ;
  assign n359 = x[67] & n330 ;
  assign n446 = x[68] & n390 ;
  assign n14068 = n359 | n446 ;
  assign n14069 = x[69] & n322 ;
  assign n14070 = n14068 | n14069 ;
  assign n14071 = n6382 | n14070 ;
  assign n28544 = ~n14071 ;
  assign n14072 = x[26] & n28544 ;
  assign n14073 = n28342 & n14071 ;
  assign n14074 = n14072 | n14073 ;
  assign n14126 = n14067 | n14074 ;
  assign n14075 = n14067 & n14074 ;
  assign n14123 = n14109 & n14121 ;
  assign n14124 = n14116 & n14118 ;
  assign n14125 = n14123 | n14124 ;
  assign n14127 = n14125 & n14126 ;
  assign n14129 = n14075 | n14127 ;
  assign n28545 = ~n14129 ;
  assign n14130 = n14126 & n28545 ;
  assign n28546 = ~n14075 ;
  assign n14128 = n28546 & n14126 ;
  assign n28547 = ~n14128 ;
  assign n14964 = n14125 & n28547 ;
  assign n14965 = n14130 | n14964 ;
  assign n5334 = n3701 & n5302 ;
  assign n5248 = x[70] & n5240 ;
  assign n6273 = x[71] & n6179 ;
  assign n14966 = n5248 | n6273 ;
  assign n14967 = x[72] & n5238 ;
  assign n14968 = n14966 | n14967 ;
  assign n14969 = n5334 | n14968 ;
  assign n28548 = ~n14969 ;
  assign n14970 = x[23] & n28548 ;
  assign n14971 = n28221 & n14969 ;
  assign n14972 = n14970 | n14971 ;
  assign n14973 = n14965 | n14972 ;
  assign n14974 = n14965 & n14972 ;
  assign n28549 = ~n14974 ;
  assign n15751 = n14973 & n28549 ;
  assign n28550 = ~n15068 ;
  assign n15753 = n28550 & n15751 ;
  assign n28551 = ~n15751 ;
  assign n15995 = n15068 & n28551 ;
  assign n15996 = n15753 | n15995 ;
  assign n15997 = n15994 & n15996 ;
  assign n16135 = n15994 | n15996 ;
  assign n28552 = ~n15997 ;
  assign n16136 = n28552 & n16135 ;
  assign n16137 = n16134 & n16136 ;
  assign n16907 = n16134 | n16136 ;
  assign n28553 = ~n16137 ;
  assign n16908 = n28553 & n16907 ;
  assign n16909 = n16906 & n16908 ;
  assign n17766 = n16906 | n16908 ;
  assign n28554 = ~n16909 ;
  assign n17767 = n28554 & n17766 ;
  assign n28555 = ~n17097 ;
  assign n17768 = n28555 & n17767 ;
  assign n28556 = ~n17767 ;
  assign n17936 = n17097 & n28556 ;
  assign n17937 = n17768 | n17936 ;
  assign n17938 = n17933 | n17937 ;
  assign n17939 = n17933 & n17937 ;
  assign n28557 = ~n17939 ;
  assign n17940 = n17938 & n28557 ;
  assign n19064 = n17949 & n17952 ;
  assign n19119 = n17965 | n19118 ;
  assign n19120 = n19065 & n19119 ;
  assign n19121 = n19064 | n19120 ;
  assign n28558 = ~n19121 ;
  assign n19122 = n17940 & n28558 ;
  assign n28559 = ~n17940 ;
  assign n19170 = n28559 & n19121 ;
  assign n19171 = n19122 | n19170 ;
  assign n12708 = n1293 & n12695 ;
  assign n12647 = x[82] & n12633 ;
  assign n14365 = x[83] & n13533 ;
  assign n19172 = n12647 | n14365 ;
  assign n19173 = x[84] & n12631 ;
  assign n19174 = n19172 | n19173 ;
  assign n19175 = n12708 | n19174 ;
  assign n28560 = ~n19175 ;
  assign n19176 = x[11] & n28560 ;
  assign n19177 = n27892 & n19175 ;
  assign n19178 = n19176 | n19177 ;
  assign n19458 = n19171 | n19178 ;
  assign n28561 = ~n16906 ;
  assign n16910 = n28561 & n16908 ;
  assign n28562 = ~n16908 ;
  assign n16911 = n16906 & n28562 ;
  assign n16912 = n16910 | n16911 ;
  assign n17098 = n16912 | n17097 ;
  assign n17099 = n16912 & n17097 ;
  assign n28563 = ~n17099 ;
  assign n17926 = n17098 & n28563 ;
  assign n28564 = ~n17933 ;
  assign n17934 = n17926 & n28564 ;
  assign n28565 = ~n17926 ;
  assign n19062 = n28565 & n17933 ;
  assign n19063 = n17934 | n19062 ;
  assign n19123 = n19063 | n19121 ;
  assign n19124 = n19063 & n19121 ;
  assign n28566 = ~n19124 ;
  assign n20322 = n19123 & n28566 ;
  assign n20323 = n19178 & n20322 ;
  assign n28567 = ~n20323 ;
  assign n20475 = n19458 & n28567 ;
  assign n28568 = ~n20475 ;
  assign n20476 = n20390 & n28568 ;
  assign n19179 = n19171 & n19178 ;
  assign n19189 = n19180 & n19187 ;
  assign n19192 = n19187 | n19191 ;
  assign n28569 = ~n19193 ;
  assign n19194 = n19192 & n28569 ;
  assign n19455 = n19205 | n19454 ;
  assign n19456 = n19194 & n19455 ;
  assign n19457 = n19189 | n19456 ;
  assign n19459 = n19457 & n19458 ;
  assign n19460 = n19179 | n19459 ;
  assign n28570 = ~n19460 ;
  assign n20477 = n19458 & n28570 ;
  assign n20478 = n20476 | n20477 ;
  assign n15325 = n1522 & n15308 ;
  assign n15257 = x[85] & n15246 ;
  assign n17291 = x[86] & n16288 ;
  assign n20479 = n15257 | n17291 ;
  assign n20480 = x[87] & n15244 ;
  assign n20481 = n20479 | n20480 ;
  assign n20482 = n15325 | n20481 ;
  assign n28571 = ~n20482 ;
  assign n20483 = x[8] & n28571 ;
  assign n20484 = n27845 & n20482 ;
  assign n20485 = n20483 | n20484 ;
  assign n28572 = ~n20485 ;
  assign n20486 = n20478 & n28572 ;
  assign n28573 = ~n20478 ;
  assign n20488 = n28573 & n20485 ;
  assign n20489 = n20486 | n20488 ;
  assign n21133 = n20498 & n20501 ;
  assign n28574 = ~n20386 ;
  assign n20387 = n19194 & n28574 ;
  assign n28575 = ~n19194 ;
  assign n20490 = n28575 & n20386 ;
  assign n20491 = n20387 | n20490 ;
  assign n20499 = n20491 | n20498 ;
  assign n20500 = n20491 & n20498 ;
  assign n28576 = ~n20500 ;
  assign n21134 = n20499 & n28576 ;
  assign n21215 = n20518 | n21214 ;
  assign n21216 = n21134 & n21215 ;
  assign n21217 = n21133 | n21216 ;
  assign n21219 = n20489 | n21217 ;
  assign n21220 = n20489 & n21217 ;
  assign n28577 = ~n21220 ;
  assign n21925 = n21219 & n28577 ;
  assign n28578 = ~n21542 ;
  assign n21926 = n28578 & n21925 ;
  assign n28579 = ~n21925 ;
  assign n21928 = n21542 & n28579 ;
  assign n21929 = n21926 | n21928 ;
  assign n28580 = ~n20810 ;
  assign n21135 = n28580 & n21134 ;
  assign n28581 = ~n21134 ;
  assign n21553 = n20810 & n28581 ;
  assign n21554 = n21135 | n21553 ;
  assign n21555 = n21552 & n21554 ;
  assign n28582 = ~n21552 ;
  assign n21558 = n28582 & n21556 ;
  assign n28583 = ~n21556 ;
  assign n22120 = n21552 & n28583 ;
  assign n22121 = n21558 | n22120 ;
  assign n22220 = n22121 & n22218 ;
  assign n22221 = n21555 | n22220 ;
  assign n28584 = ~n21929 ;
  assign n22222 = n28584 & n22221 ;
  assign n28585 = ~n22221 ;
  assign n22520 = n21929 & n28585 ;
  assign n22521 = n22222 | n22520 ;
  assign n540 = n538 & n539 ;
  assign n541 = n26068 | n540 ;
  assign n27631 = x[92] & x[93] ;
  assign n542 = x[92] | x[93] ;
  assign n28586 = ~n27631 ;
  assign n1682 = n28586 & n542 ;
  assign n28587 = ~n541 ;
  assign n1683 = n28587 & n1682 ;
  assign n28588 = ~n1682 ;
  assign n1684 = n541 & n28588 ;
  assign n1685 = n1683 | n1684 ;
  assign n19703 = n1685 & n19656 ;
  assign n19743 = x[91] & n19723 ;
  assign n19847 = x[92] & n19829 ;
  assign n22522 = n19743 | n19847 ;
  assign n22523 = x[93] & n19655 ;
  assign n22524 = n22522 | n22523 ;
  assign n22525 = n19703 | n22524 ;
  assign n28589 = ~n22525 ;
  assign n22526 = x[2] & n28589 ;
  assign n22527 = n27790 & n22525 ;
  assign n22528 = n22526 | n22527 ;
  assign n28590 = ~n22528 ;
  assign n22529 = n22521 & n28590 ;
  assign n28591 = ~n22521 ;
  assign n22531 = n28591 & n22528 ;
  assign n22532 = n22529 | n22531 ;
  assign n22934 = n22543 | n22933 ;
  assign n22935 = n22532 | n22934 ;
  assign n22936 = n22532 & n22934 ;
  assign n28592 = ~n22936 ;
  assign n158 = n22935 & n28592 ;
  assign n20487 = n20478 & n20485 ;
  assign n21221 = n20487 | n21220 ;
  assign n20391 = n19178 | n20322 ;
  assign n20392 = n20390 & n20391 ;
  assign n20393 = n20323 | n20392 ;
  assign n10554 = n1003 & n10542 ;
  assign n10493 = x[80] & n10481 ;
  assign n11922 = x[81] & n11232 ;
  assign n17913 = n10493 | n11922 ;
  assign n17914 = x[82] & n10479 ;
  assign n17915 = n17913 | n17914 ;
  assign n17916 = n10554 | n17915 ;
  assign n28593 = ~n17916 ;
  assign n17917 = x[14] & n28593 ;
  assign n17918 = n27956 & n17916 ;
  assign n17919 = n17917 | n17918 ;
  assign n8726 = n1741 & n8706 ;
  assign n8655 = x[77] & n8645 ;
  assign n9872 = x[78] & n9278 ;
  assign n16887 = n8655 | n9872 ;
  assign n16888 = x[79] & n8643 ;
  assign n16889 = n16887 | n16888 ;
  assign n16890 = n8726 | n16889 ;
  assign n28594 = ~n16890 ;
  assign n16891 = x[17] & n28594 ;
  assign n16892 = n28039 & n16890 ;
  assign n16893 = n16891 | n16892 ;
  assign n16138 = n15997 | n16137 ;
  assign n7168 = n2750 & n7162 ;
  assign n7106 = x[74] & n7100 ;
  assign n7679 = x[75] & n7647 ;
  assign n15978 = n7106 | n7679 ;
  assign n15979 = x[76] & n7098 ;
  assign n15980 = n15978 | n15979 ;
  assign n15981 = n7168 | n15980 ;
  assign n28595 = ~n15981 ;
  assign n15982 = x[20] & n28595 ;
  assign n15983 = n28114 & n15981 ;
  assign n15984 = n15982 | n15983 ;
  assign n5340 = n3733 & n5302 ;
  assign n5242 = x[71] & n5240 ;
  assign n6223 = x[72] & n6179 ;
  assign n14956 = n5242 | n6223 ;
  assign n14957 = x[73] & n5238 ;
  assign n14958 = n14956 | n14957 ;
  assign n14959 = n5340 | n14958 ;
  assign n28596 = ~n14959 ;
  assign n14960 = x[23] & n28596 ;
  assign n14961 = n28221 & n14959 ;
  assign n14962 = n14960 | n14961 ;
  assign n5977 = n452 & n5976 ;
  assign n336 = x[68] & n330 ;
  assign n425 = x[69] & n390 ;
  assign n14056 = n336 | n425 ;
  assign n14057 = x[70] & n322 ;
  assign n14058 = n14056 | n14057 ;
  assign n14059 = n5977 | n14058 ;
  assign n28597 = ~n14059 ;
  assign n14060 = x[26] & n28597 ;
  assign n14061 = n28342 & n14059 ;
  assign n14062 = n14060 | n14061 ;
  assign n27659 = x[29] & x[30] ;
  assign n648 = x[29] | x[30] ;
  assign n28598 = ~n27659 ;
  assign n649 = n28598 & n648 ;
  assign n12401 = x[64] & n649 ;
  assign n13318 = n12401 & n28543 ;
  assign n28599 = ~n12401 ;
  assign n13319 = n28599 & n13317 ;
  assign n13320 = n13318 | n13319 ;
  assign n6499 = n4632 & n6494 ;
  assign n4569 = x[65] & n4514 ;
  assign n4627 = x[66] & n4572 ;
  assign n13321 = n4569 | n4627 ;
  assign n13322 = x[67] & n4504 ;
  assign n13323 = n13321 | n13322 ;
  assign n13324 = n6499 | n13323 ;
  assign n28600 = ~n13324 ;
  assign n13325 = x[29] & n28600 ;
  assign n13326 = n28483 & n13324 ;
  assign n13327 = n13325 | n13326 ;
  assign n28601 = ~n13327 ;
  assign n13328 = n13320 & n28601 ;
  assign n28602 = ~n13320 ;
  assign n14063 = n28602 & n13327 ;
  assign n14064 = n13328 | n14063 ;
  assign n28603 = ~n14062 ;
  assign n14065 = n28603 & n14064 ;
  assign n28604 = ~n14064 ;
  assign n14131 = n14062 & n28604 ;
  assign n14132 = n14065 | n14131 ;
  assign n28605 = ~n14132 ;
  assign n15069 = n14129 & n28605 ;
  assign n15072 = n28545 & n14132 ;
  assign n15073 = n15069 | n15072 ;
  assign n15074 = n14962 & n15073 ;
  assign n14133 = n14129 | n14132 ;
  assign n14134 = n14129 & n14132 ;
  assign n28606 = ~n14134 ;
  assign n14955 = n14133 & n28606 ;
  assign n15075 = n14955 | n14962 ;
  assign n28607 = ~n15074 ;
  assign n15076 = n28607 & n15075 ;
  assign n15749 = n15064 & n15065 ;
  assign n15750 = n14984 | n15749 ;
  assign n15752 = n15750 & n15751 ;
  assign n15754 = n14974 | n15752 ;
  assign n28608 = ~n15754 ;
  assign n15755 = n15076 & n28608 ;
  assign n28609 = ~n15076 ;
  assign n15985 = n28609 & n15754 ;
  assign n15986 = n15755 | n15985 ;
  assign n15987 = n15984 & n15986 ;
  assign n16139 = n15984 | n15986 ;
  assign n28610 = ~n15987 ;
  assign n16436 = n28610 & n16139 ;
  assign n28611 = ~n16138 ;
  assign n16438 = n28611 & n16436 ;
  assign n28612 = ~n16436 ;
  assign n16894 = n16138 & n28612 ;
  assign n16895 = n16438 | n16894 ;
  assign n28613 = ~n16893 ;
  assign n16897 = n28613 & n16895 ;
  assign n28614 = ~n16895 ;
  assign n17764 = n16893 & n28614 ;
  assign n17765 = n16897 | n17764 ;
  assign n17792 = n16926 | n17791 ;
  assign n17793 = n17767 & n17792 ;
  assign n17794 = n16909 | n17793 ;
  assign n17796 = n17765 | n17794 ;
  assign n17797 = n17765 & n17794 ;
  assign n28615 = ~n17797 ;
  assign n17922 = n17796 & n28615 ;
  assign n28616 = ~n17919 ;
  assign n17923 = n28616 & n17922 ;
  assign n28617 = ~n17922 ;
  assign n17924 = n17919 & n28617 ;
  assign n17925 = n17923 | n17924 ;
  assign n17935 = n17926 & n17933 ;
  assign n18170 = n17951 | n18169 ;
  assign n18171 = n17940 & n18170 ;
  assign n18172 = n17935 | n18171 ;
  assign n18173 = n17925 | n18172 ;
  assign n18174 = n17925 & n18172 ;
  assign n28618 = ~n18174 ;
  assign n19160 = n18173 & n28618 ;
  assign n12709 = n1239 & n12695 ;
  assign n12691 = x[83] & n12633 ;
  assign n14366 = x[84] & n13533 ;
  assign n19161 = n12691 | n14366 ;
  assign n19162 = x[85] & n12631 ;
  assign n19163 = n19161 | n19162 ;
  assign n19164 = n12709 | n19163 ;
  assign n28619 = ~n19164 ;
  assign n19165 = x[11] & n28619 ;
  assign n19166 = n27892 & n19164 ;
  assign n19167 = n19165 | n19166 ;
  assign n28620 = ~n19167 ;
  assign n19168 = n19160 & n28620 ;
  assign n28621 = ~n19160 ;
  assign n20394 = n28621 & n19167 ;
  assign n20395 = n19168 | n20394 ;
  assign n20396 = n20393 | n20395 ;
  assign n20397 = n20393 & n20395 ;
  assign n28622 = ~n20397 ;
  assign n20466 = n20396 & n28622 ;
  assign n15363 = n1720 & n15308 ;
  assign n15291 = x[86] & n15246 ;
  assign n17289 = x[87] & n16288 ;
  assign n20467 = n15291 | n17289 ;
  assign n20468 = x[88] & n15244 ;
  assign n20469 = n20467 | n20468 ;
  assign n20470 = n15363 | n20469 ;
  assign n28623 = ~n20470 ;
  assign n20471 = x[8] & n28623 ;
  assign n20472 = n27845 & n20470 ;
  assign n20473 = n20471 | n20472 ;
  assign n20474 = n20466 & n20473 ;
  assign n20816 = n20466 | n20473 ;
  assign n28624 = ~n20474 ;
  assign n21222 = n28624 & n20816 ;
  assign n21223 = n21221 & n21222 ;
  assign n21523 = n21221 | n21222 ;
  assign n28625 = ~n21223 ;
  assign n21524 = n28625 & n21523 ;
  assign n18408 = n2046 & n18392 ;
  assign n18340 = x[89] & n18329 ;
  assign n18529 = x[90] & n18514 ;
  assign n21525 = n18340 | n18529 ;
  assign n21526 = x[91] & n18327 ;
  assign n21527 = n21525 | n21526 ;
  assign n21528 = n18408 | n21527 ;
  assign n28626 = ~n21528 ;
  assign n21529 = x[5] & n28626 ;
  assign n21530 = n27813 & n21528 ;
  assign n21531 = n21529 | n21530 ;
  assign n28627 = ~n21531 ;
  assign n21532 = n21524 & n28627 ;
  assign n28628 = ~n21524 ;
  assign n22118 = n28628 & n21531 ;
  assign n22119 = n21532 | n22118 ;
  assign n28629 = ~n21217 ;
  assign n21218 = n20489 & n28629 ;
  assign n28630 = ~n20489 ;
  assign n21543 = n28630 & n21217 ;
  assign n21544 = n21218 | n21543 ;
  assign n21545 = n21542 & n21544 ;
  assign n21927 = n21542 & n21925 ;
  assign n22223 = n21542 | n21925 ;
  assign n28631 = ~n21927 ;
  assign n22224 = n28631 & n22223 ;
  assign n22225 = n22221 & n22224 ;
  assign n22226 = n21545 | n22225 ;
  assign n22227 = n22119 | n22226 ;
  assign n22228 = n22119 & n22226 ;
  assign n28632 = ~n22228 ;
  assign n22508 = n22227 & n28632 ;
  assign n543 = n541 & n542 ;
  assign n544 = n27631 | n543 ;
  assign n25940 = x[93] & x[94] ;
  assign n545 = x[93] | x[94] ;
  assign n28633 = ~n25940 ;
  assign n2407 = n28633 & n545 ;
  assign n2408 = n544 & n2407 ;
  assign n2409 = n544 | n2407 ;
  assign n28634 = ~n2408 ;
  assign n2410 = n28634 & n2409 ;
  assign n19712 = n2410 & n19656 ;
  assign n19747 = x[92] & n19723 ;
  assign n19861 = x[93] & n19829 ;
  assign n22509 = n19747 | n19861 ;
  assign n22510 = x[94] & n19655 ;
  assign n22511 = n22509 | n22510 ;
  assign n22512 = n19712 | n22511 ;
  assign n28635 = ~n22512 ;
  assign n22513 = x[2] & n28635 ;
  assign n22514 = n27790 & n22512 ;
  assign n22515 = n22513 | n22514 ;
  assign n28636 = ~n22515 ;
  assign n22516 = n22508 & n28636 ;
  assign n28637 = ~n22508 ;
  assign n22518 = n28637 & n22515 ;
  assign n22519 = n22516 | n22518 ;
  assign n22530 = n22521 & n22528 ;
  assign n22937 = n22530 | n22936 ;
  assign n22938 = n22519 & n22937 ;
  assign n27666 = n22519 | n22937 ;
  assign n28638 = ~n22938 ;
  assign n159 = n28638 & n27666 ;
  assign n21533 = n21524 & n21531 ;
  assign n21534 = n21524 | n21531 ;
  assign n28639 = ~n21533 ;
  assign n21535 = n28639 & n21534 ;
  assign n28640 = ~n21567 ;
  assign n21572 = n28640 & n21571 ;
  assign n28641 = ~n21571 ;
  assign n21574 = n21567 & n28641 ;
  assign n21575 = n21572 | n21574 ;
  assign n21921 = n21575 & n21920 ;
  assign n21922 = n21570 | n21921 ;
  assign n21923 = n21560 & n21922 ;
  assign n21924 = n21555 | n21923 ;
  assign n21930 = n21924 & n21929 ;
  assign n21931 = n21545 | n21930 ;
  assign n21932 = n21535 & n21931 ;
  assign n21933 = n21533 | n21932 ;
  assign n15326 = n1453 & n15308 ;
  assign n15294 = x[87] & n15246 ;
  assign n17294 = x[88] & n16288 ;
  assign n20452 = n15294 | n17294 ;
  assign n20453 = x[89] & n15244 ;
  assign n20454 = n20452 | n20453 ;
  assign n20455 = n15326 | n20454 ;
  assign n28642 = ~n20455 ;
  assign n20456 = x[8] & n28642 ;
  assign n20457 = n27845 & n20455 ;
  assign n20458 = n20456 | n20457 ;
  assign n19169 = n19160 & n19167 ;
  assign n16896 = n16893 & n16895 ;
  assign n16898 = n16893 | n16895 ;
  assign n28643 = ~n16896 ;
  assign n16899 = n28643 & n16898 ;
  assign n28644 = ~n17794 ;
  assign n17795 = n16899 & n28644 ;
  assign n28645 = ~n16899 ;
  assign n17911 = n28645 & n17794 ;
  assign n17912 = n17795 | n17911 ;
  assign n17920 = n17912 | n17919 ;
  assign n17921 = n17912 & n17919 ;
  assign n28646 = ~n17921 ;
  assign n19060 = n17920 & n28646 ;
  assign n28647 = ~n18172 ;
  assign n19061 = n28647 & n19060 ;
  assign n28648 = ~n19060 ;
  assign n19461 = n18172 & n28648 ;
  assign n19462 = n19061 | n19461 ;
  assign n19463 = n19167 | n19462 ;
  assign n19464 = n19167 & n19462 ;
  assign n28649 = ~n19464 ;
  assign n19465 = n19463 & n28649 ;
  assign n19466 = n19460 & n19465 ;
  assign n19467 = n19169 | n19466 ;
  assign n17100 = n16909 | n17099 ;
  assign n17101 = n16899 & n17100 ;
  assign n17102 = n16896 | n17101 ;
  assign n8729 = n1270 & n8706 ;
  assign n8676 = x[78] & n8645 ;
  assign n9884 = x[79] & n9278 ;
  assign n16872 = n8676 | n9884 ;
  assign n16873 = x[80] & n8643 ;
  assign n16874 = n16872 | n16873 ;
  assign n16875 = n8729 | n16874 ;
  assign n28650 = ~n16875 ;
  assign n16876 = x[17] & n28650 ;
  assign n16877 = n28039 & n16875 ;
  assign n16878 = n16876 | n16877 ;
  assign n14066 = n14062 & n14064 ;
  assign n14135 = n14066 | n14134 ;
  assign n4797 = n452 & n4790 ;
  assign n333 = x[69] & n330 ;
  assign n445 = x[70] & n390 ;
  assign n14045 = n333 | n445 ;
  assign n14046 = x[71] & n322 ;
  assign n14047 = n14045 | n14046 ;
  assign n14048 = n4797 | n14047 ;
  assign n28651 = ~n14048 ;
  assign n14049 = x[26] & n28651 ;
  assign n14050 = n28342 & n14048 ;
  assign n14051 = n14049 | n14050 ;
  assign n13329 = n13320 & n13327 ;
  assign n13330 = n12401 & n13317 ;
  assign n13331 = n13329 | n13330 ;
  assign n6416 = n4632 & n6408 ;
  assign n4543 = x[66] & n4514 ;
  assign n4628 = x[67] & n4572 ;
  assign n13332 = n4543 | n4628 ;
  assign n13333 = x[68] & n4504 ;
  assign n13334 = n13332 | n13333 ;
  assign n13335 = n6416 | n13334 ;
  assign n28652 = ~n13335 ;
  assign n13336 = x[29] & n28652 ;
  assign n13337 = n28483 & n13335 ;
  assign n13338 = n13336 | n13337 ;
  assign n12402 = x[32] & n28599 ;
  assign n27661 = x[31] & x[32] ;
  assign n650 = x[31] | x[32] ;
  assign n28653 = ~n27661 ;
  assign n651 = n28653 & n650 ;
  assign n779 = n649 & n651 ;
  assign n6439 = n779 & n6437 ;
  assign n28654 = ~n651 ;
  assign n652 = n649 & n28654 ;
  assign n12403 = x[65] & n652 ;
  assign n27662 = x[30] & x[31] ;
  assign n660 = x[30] | x[31] ;
  assign n28655 = ~n27662 ;
  assign n661 = n28655 & n660 ;
  assign n28656 = ~n649 ;
  assign n720 = n28656 & n661 ;
  assign n12404 = x[64] & n720 ;
  assign n12405 = n12403 | n12404 ;
  assign n12406 = n6439 | n12405 ;
  assign n28657 = ~n12406 ;
  assign n12407 = x[32] & n28657 ;
  assign n28658 = ~x[32] ;
  assign n12408 = n28658 & n12406 ;
  assign n12409 = n12407 | n12408 ;
  assign n28659 = ~n12409 ;
  assign n12410 = n12402 & n28659 ;
  assign n28660 = ~n12402 ;
  assign n13339 = n28660 & n12409 ;
  assign n13340 = n12410 | n13339 ;
  assign n28661 = ~n13338 ;
  assign n13341 = n28661 & n13340 ;
  assign n28662 = ~n13340 ;
  assign n13342 = n13338 & n28662 ;
  assign n13343 = n13341 | n13342 ;
  assign n28663 = ~n13343 ;
  assign n13344 = n13331 & n28663 ;
  assign n28664 = ~n13331 ;
  assign n14052 = n28664 & n13343 ;
  assign n14053 = n13344 | n14052 ;
  assign n14054 = n14051 | n14053 ;
  assign n14055 = n14051 & n14053 ;
  assign n28665 = ~n14055 ;
  assign n14136 = n14054 & n28665 ;
  assign n14137 = n14135 & n14136 ;
  assign n14941 = n14135 | n14136 ;
  assign n28666 = ~n14137 ;
  assign n14942 = n28666 & n14941 ;
  assign n5309 = n2722 & n5302 ;
  assign n5290 = x[72] & n5240 ;
  assign n6224 = x[73] & n6179 ;
  assign n14943 = n5290 | n6224 ;
  assign n14944 = x[74] & n5238 ;
  assign n14945 = n14943 | n14944 ;
  assign n14946 = n5309 | n14945 ;
  assign n28667 = ~n14946 ;
  assign n14947 = x[23] & n28667 ;
  assign n14948 = n28221 & n14946 ;
  assign n14949 = n14947 | n14948 ;
  assign n28668 = ~n14949 ;
  assign n14952 = n14942 & n28668 ;
  assign n28669 = ~n14942 ;
  assign n14953 = n28669 & n14949 ;
  assign n14954 = n14952 | n14953 ;
  assign n14963 = n14955 & n14962 ;
  assign n15070 = n14973 & n15068 ;
  assign n15071 = n14974 | n15070 ;
  assign n15077 = n15071 & n15076 ;
  assign n15078 = n14963 | n15077 ;
  assign n15079 = n14954 | n15078 ;
  assign n15080 = n14954 & n15078 ;
  assign n28670 = ~n15080 ;
  assign n15963 = n15079 & n28670 ;
  assign n7189 = n1775 & n7162 ;
  assign n7141 = x[75] & n7100 ;
  assign n7680 = x[76] & n7647 ;
  assign n15964 = n7141 | n7680 ;
  assign n15965 = x[77] & n7098 ;
  assign n15966 = n15964 | n15965 ;
  assign n15967 = n7189 | n15966 ;
  assign n28671 = ~n15967 ;
  assign n15968 = x[20] & n28671 ;
  assign n15969 = n28114 & n15967 ;
  assign n15970 = n15968 | n15969 ;
  assign n28672 = ~n15970 ;
  assign n15971 = n15963 & n28672 ;
  assign n28673 = ~n15963 ;
  assign n16421 = n28673 & n15970 ;
  assign n16422 = n15971 | n16421 ;
  assign n16430 = n16128 & n16428 ;
  assign n16431 = n16127 | n16430 ;
  assign n16432 = n16423 & n16431 ;
  assign n16433 = n16008 | n16432 ;
  assign n16434 = n16135 & n16433 ;
  assign n16435 = n15997 | n16434 ;
  assign n16437 = n16435 & n16436 ;
  assign n16439 = n15987 | n16437 ;
  assign n16441 = n16422 | n16439 ;
  assign n16442 = n16422 & n16439 ;
  assign n28674 = ~n16442 ;
  assign n16882 = n16441 & n28674 ;
  assign n16884 = n16878 & n16882 ;
  assign n17761 = n16878 | n16882 ;
  assign n28675 = ~n16884 ;
  assign n17762 = n28675 & n17761 ;
  assign n28676 = ~n17102 ;
  assign n17763 = n28676 & n17762 ;
  assign n28677 = ~n17762 ;
  assign n17899 = n17102 & n28677 ;
  assign n17900 = n17763 | n17899 ;
  assign n10599 = n1057 & n10542 ;
  assign n10494 = x[81] & n10481 ;
  assign n11914 = x[82] & n11232 ;
  assign n17901 = n10494 | n11914 ;
  assign n17902 = x[83] & n10479 ;
  assign n17903 = n17901 | n17902 ;
  assign n17904 = n10599 | n17903 ;
  assign n28678 = ~n17904 ;
  assign n17905 = x[14] & n28678 ;
  assign n17906 = n27956 & n17904 ;
  assign n17907 = n17905 | n17906 ;
  assign n17908 = n17900 | n17907 ;
  assign n17909 = n17900 & n17907 ;
  assign n28679 = ~n17909 ;
  assign n17910 = n17908 & n28679 ;
  assign n19059 = n17919 & n17922 ;
  assign n19125 = n17939 | n19124 ;
  assign n19126 = n19060 & n19125 ;
  assign n19127 = n19059 | n19126 ;
  assign n28680 = ~n19127 ;
  assign n19128 = n17910 & n28680 ;
  assign n28681 = ~n17910 ;
  assign n19144 = n28681 & n19127 ;
  assign n19145 = n19128 | n19144 ;
  assign n12711 = n1213 & n12695 ;
  assign n12683 = x[84] & n12633 ;
  assign n14369 = x[85] & n13533 ;
  assign n19146 = n12683 | n14369 ;
  assign n19147 = x[86] & n12631 ;
  assign n19148 = n19146 | n19147 ;
  assign n19149 = n12711 | n19148 ;
  assign n28682 = ~n19149 ;
  assign n19150 = x[11] & n28682 ;
  assign n19151 = n27892 & n19149 ;
  assign n19152 = n19150 | n19151 ;
  assign n19153 = n19145 | n19152 ;
  assign n19154 = n19145 & n19152 ;
  assign n28683 = ~n19154 ;
  assign n20320 = n19153 & n28683 ;
  assign n28684 = ~n19467 ;
  assign n20321 = n28684 & n20320 ;
  assign n28685 = ~n20320 ;
  assign n20461 = n19467 & n28685 ;
  assign n20462 = n20321 | n20461 ;
  assign n20463 = n20458 | n20462 ;
  assign n20464 = n20458 & n20462 ;
  assign n28686 = ~n20464 ;
  assign n20465 = n20463 & n28686 ;
  assign n21224 = n20474 | n21223 ;
  assign n28687 = ~n21224 ;
  assign n21225 = n20465 & n28687 ;
  assign n28688 = ~n20465 ;
  assign n21508 = n28688 & n21224 ;
  assign n21509 = n21225 | n21508 ;
  assign n18439 = n1841 & n18392 ;
  assign n18343 = x[90] & n18329 ;
  assign n18553 = x[91] & n18514 ;
  assign n21510 = n18343 | n18553 ;
  assign n21511 = x[92] & n18327 ;
  assign n21512 = n21510 | n21511 ;
  assign n21513 = n18439 | n21512 ;
  assign n28689 = ~n21513 ;
  assign n21514 = x[5] & n28689 ;
  assign n21515 = n27813 & n21513 ;
  assign n21516 = n21514 | n21515 ;
  assign n21517 = n21509 | n21516 ;
  assign n21518 = n21509 & n21516 ;
  assign n28690 = ~n21518 ;
  assign n22116 = n21517 & n28690 ;
  assign n28691 = ~n21933 ;
  assign n22117 = n28691 & n22116 ;
  assign n28692 = ~n22116 ;
  assign n22496 = n21933 & n28692 ;
  assign n22497 = n22117 | n22496 ;
  assign n546 = n544 & n545 ;
  assign n547 = n25940 | n546 ;
  assign n27630 = x[94] & x[95] ;
  assign n548 = x[94] | x[95] ;
  assign n28693 = ~n27630 ;
  assign n2149 = n28693 & n548 ;
  assign n2150 = n547 | n2149 ;
  assign n2151 = n547 & n2149 ;
  assign n28694 = ~n2151 ;
  assign n2152 = n2150 & n28694 ;
  assign n19699 = n2152 & n19656 ;
  assign n19746 = x[93] & n19723 ;
  assign n19845 = x[94] & n19829 ;
  assign n22498 = n19746 | n19845 ;
  assign n22499 = x[95] & n19655 ;
  assign n22500 = n22498 | n22499 ;
  assign n22501 = n19699 | n22500 ;
  assign n28695 = ~n22501 ;
  assign n22502 = x[2] & n28695 ;
  assign n22503 = n27790 & n22501 ;
  assign n22504 = n22502 | n22503 ;
  assign n22505 = n22497 | n22504 ;
  assign n22506 = n22497 & n22504 ;
  assign n28696 = ~n22506 ;
  assign n22507 = n22505 & n28696 ;
  assign n22517 = n22508 & n22515 ;
  assign n22939 = n22517 | n22938 ;
  assign n22940 = n22507 | n22939 ;
  assign n22941 = n22507 & n22939 ;
  assign n28697 = ~n22941 ;
  assign n160 = n22940 & n28697 ;
  assign n22942 = n22506 | n22941 ;
  assign n18175 = n17921 | n18174 ;
  assign n18176 = n17910 & n18175 ;
  assign n19155 = n17910 | n18175 ;
  assign n28698 = ~n18176 ;
  assign n19156 = n28698 & n19155 ;
  assign n28699 = ~n19152 ;
  assign n19157 = n28699 & n19156 ;
  assign n28700 = ~n19156 ;
  assign n19158 = n19152 & n28700 ;
  assign n19159 = n19157 | n19158 ;
  assign n19468 = n19159 | n19467 ;
  assign n19469 = n19159 & n19467 ;
  assign n28701 = ~n19469 ;
  assign n20451 = n19468 & n28701 ;
  assign n28702 = ~n20458 ;
  assign n20459 = n20451 & n28702 ;
  assign n28703 = ~n20451 ;
  assign n21131 = n28703 & n20458 ;
  assign n21132 = n20459 | n21131 ;
  assign n21226 = n21132 | n21224 ;
  assign n21227 = n21132 & n21224 ;
  assign n28704 = ~n21227 ;
  assign n21519 = n21226 & n28704 ;
  assign n28705 = ~n21516 ;
  assign n21520 = n28705 & n21519 ;
  assign n28706 = ~n21519 ;
  assign n21521 = n21516 & n28706 ;
  assign n21522 = n21520 | n21521 ;
  assign n21934 = n21522 & n21933 ;
  assign n21935 = n21518 | n21934 ;
  assign n15329 = n1482 & n15308 ;
  assign n15279 = x[88] & n15246 ;
  assign n17290 = x[89] & n16288 ;
  assign n20438 = n15279 | n17290 ;
  assign n20439 = x[90] & n15244 ;
  assign n20440 = n20438 | n20439 ;
  assign n20441 = n15329 | n20440 ;
  assign n28707 = ~n20441 ;
  assign n20442 = x[8] & n28707 ;
  assign n20443 = n27845 & n20441 ;
  assign n20444 = n20442 | n20443 ;
  assign n19470 = n19154 | n19469 ;
  assign n19129 = n17910 & n19127 ;
  assign n19130 = n17909 | n19129 ;
  assign n8712 = n1029 & n8706 ;
  assign n8682 = x[79] & n8645 ;
  assign n9892 = x[80] & n9278 ;
  assign n16859 = n8682 | n9892 ;
  assign n16860 = x[81] & n8643 ;
  assign n16861 = n16859 | n16860 ;
  assign n16862 = n8712 | n16861 ;
  assign n28708 = ~n16862 ;
  assign n16863 = x[17] & n28708 ;
  assign n16864 = n28039 & n16862 ;
  assign n16865 = n16863 | n16864 ;
  assign n14950 = n14942 | n14949 ;
  assign n14951 = n14942 & n14949 ;
  assign n28709 = ~n14951 ;
  assign n15746 = n14950 & n28709 ;
  assign n28710 = ~n15078 ;
  assign n15747 = n28710 & n15746 ;
  assign n28711 = ~n15746 ;
  assign n15973 = n15078 & n28711 ;
  assign n15974 = n15747 | n15973 ;
  assign n15976 = n15970 & n15974 ;
  assign n16443 = n15976 | n16442 ;
  assign n15081 = n14951 | n15080 ;
  assign n13345 = n13331 & n13343 ;
  assign n13346 = n13338 & n13340 ;
  assign n13347 = n13345 | n13346 ;
  assign n12411 = n12402 & n12409 ;
  assign n6467 = n779 & n6466 ;
  assign n662 = n28656 & n651 ;
  assign n28712 = ~n661 ;
  assign n663 = n28712 & n662 ;
  assign n685 = x[64] & n663 ;
  assign n773 = x[65] & n720 ;
  assign n12412 = n685 | n773 ;
  assign n12413 = x[66] & n652 ;
  assign n12414 = n12412 | n12413 ;
  assign n12415 = n6467 | n12414 ;
  assign n28713 = ~n12415 ;
  assign n12416 = x[32] & n28713 ;
  assign n12417 = n28658 & n12415 ;
  assign n12418 = n12416 | n12417 ;
  assign n12419 = n12411 | n12418 ;
  assign n12420 = n12411 & n12418 ;
  assign n28714 = ~n12420 ;
  assign n13289 = n12419 & n28714 ;
  assign n6387 = n4632 & n6379 ;
  assign n4567 = x[67] & n4514 ;
  assign n4576 = x[68] & n4572 ;
  assign n13290 = n4567 | n4576 ;
  assign n13291 = x[69] & n4504 ;
  assign n13292 = n13290 | n13291 ;
  assign n13293 = n6387 | n13292 ;
  assign n28715 = ~n13293 ;
  assign n13294 = x[29] & n28715 ;
  assign n13295 = n28483 & n13293 ;
  assign n13296 = n13294 | n13295 ;
  assign n13297 = n13289 & n13296 ;
  assign n13348 = n13289 | n13296 ;
  assign n28716 = ~n13297 ;
  assign n13350 = n28716 & n13348 ;
  assign n28717 = ~n13350 ;
  assign n14030 = n13347 & n28717 ;
  assign n13349 = n13347 & n13348 ;
  assign n13351 = n13297 | n13349 ;
  assign n28718 = ~n13351 ;
  assign n14031 = n13348 & n28718 ;
  assign n14032 = n14030 | n14031 ;
  assign n3703 = n452 & n3701 ;
  assign n374 = x[70] & n330 ;
  assign n429 = x[71] & n390 ;
  assign n14033 = n374 | n429 ;
  assign n14034 = x[72] & n322 ;
  assign n14035 = n14033 | n14034 ;
  assign n14036 = n3703 | n14035 ;
  assign n28719 = ~n14036 ;
  assign n14037 = x[26] & n28719 ;
  assign n14038 = n28342 & n14036 ;
  assign n14039 = n14037 | n14038 ;
  assign n28720 = ~n14039 ;
  assign n14042 = n14032 & n28720 ;
  assign n28721 = ~n14032 ;
  assign n14043 = n28721 & n14039 ;
  assign n14044 = n14042 | n14043 ;
  assign n14138 = n14055 | n14137 ;
  assign n14139 = n14044 | n14138 ;
  assign n14140 = n14044 & n14138 ;
  assign n28722 = ~n14140 ;
  assign n14932 = n14139 & n28722 ;
  assign n5311 = n3289 & n5302 ;
  assign n5244 = x[73] & n5240 ;
  assign n6225 = x[74] & n6179 ;
  assign n14933 = n5244 | n6225 ;
  assign n14934 = x[75] & n5238 ;
  assign n14935 = n14933 | n14934 ;
  assign n14936 = n5311 | n14935 ;
  assign n28723 = ~n14936 ;
  assign n14937 = x[23] & n28723 ;
  assign n14938 = n28221 & n14936 ;
  assign n14939 = n14937 | n14938 ;
  assign n14940 = n14932 & n14939 ;
  assign n14040 = n14032 | n14039 ;
  assign n14041 = n14032 & n14039 ;
  assign n28724 = ~n14041 ;
  assign n14704 = n14040 & n28724 ;
  assign n28725 = ~n14138 ;
  assign n14705 = n28725 & n14704 ;
  assign n28726 = ~n14704 ;
  assign n15743 = n14138 & n28726 ;
  assign n15744 = n14705 | n15743 ;
  assign n15760 = n14939 | n15744 ;
  assign n28727 = ~n14940 ;
  assign n15950 = n28727 & n15760 ;
  assign n28728 = ~n15950 ;
  assign n15951 = n15081 & n28728 ;
  assign n15745 = n14939 & n15744 ;
  assign n15756 = n15075 & n15754 ;
  assign n15757 = n15074 | n15756 ;
  assign n15758 = n15746 & n15757 ;
  assign n15759 = n14951 | n15758 ;
  assign n15761 = n15759 & n15760 ;
  assign n15762 = n15745 | n15761 ;
  assign n28729 = ~n15762 ;
  assign n15952 = n15760 & n28729 ;
  assign n15953 = n15951 | n15952 ;
  assign n7169 = n2084 & n7162 ;
  assign n7107 = x[76] & n7100 ;
  assign n7720 = x[77] & n7647 ;
  assign n15954 = n7107 | n7720 ;
  assign n15955 = x[78] & n7098 ;
  assign n15956 = n15954 | n15955 ;
  assign n15957 = n7169 | n15956 ;
  assign n28730 = ~n15957 ;
  assign n15958 = x[20] & n28730 ;
  assign n15959 = n28114 & n15957 ;
  assign n15960 = n15958 | n15959 ;
  assign n28731 = ~n15960 ;
  assign n15961 = n15953 & n28731 ;
  assign n28732 = ~n15953 ;
  assign n16444 = n28732 & n15960 ;
  assign n16445 = n15961 | n16444 ;
  assign n16446 = n16443 & n16445 ;
  assign n16866 = n16443 | n16445 ;
  assign n28733 = ~n16446 ;
  assign n16867 = n28733 & n16866 ;
  assign n16868 = n16865 & n16867 ;
  assign n16870 = n16865 | n16867 ;
  assign n28734 = ~n16868 ;
  assign n16871 = n28734 & n16870 ;
  assign n15975 = n15970 | n15974 ;
  assign n28735 = ~n15976 ;
  assign n15977 = n15975 & n28735 ;
  assign n28736 = ~n16439 ;
  assign n16440 = n15977 & n28736 ;
  assign n28737 = ~n15977 ;
  assign n16879 = n28737 & n16439 ;
  assign n16880 = n16440 | n16879 ;
  assign n16881 = n16878 & n16880 ;
  assign n17798 = n16896 | n17797 ;
  assign n17799 = n17762 & n17798 ;
  assign n17800 = n16881 | n17799 ;
  assign n28738 = ~n17800 ;
  assign n17801 = n16871 & n28738 ;
  assign n28739 = ~n16871 ;
  assign n17889 = n28739 & n17800 ;
  assign n17890 = n17801 | n17889 ;
  assign n10572 = n1293 & n10542 ;
  assign n10522 = x[82] & n10481 ;
  assign n11891 = x[83] & n11232 ;
  assign n17891 = n10522 | n11891 ;
  assign n17892 = x[84] & n10479 ;
  assign n17893 = n17891 | n17892 ;
  assign n17894 = n10572 | n17893 ;
  assign n28740 = ~n17894 ;
  assign n17895 = x[14] & n28740 ;
  assign n17896 = n27956 & n17894 ;
  assign n17897 = n17895 | n17896 ;
  assign n17898 = n17890 & n17897 ;
  assign n18178 = n17890 | n17897 ;
  assign n28741 = ~n17898 ;
  assign n19131 = n28741 & n18178 ;
  assign n28742 = ~n19131 ;
  assign n19132 = n19130 & n28742 ;
  assign n18177 = n17909 | n18176 ;
  assign n18179 = n18177 & n18178 ;
  assign n18180 = n17898 | n18179 ;
  assign n28743 = ~n18180 ;
  assign n19133 = n18178 & n28743 ;
  assign n19134 = n19132 | n19133 ;
  assign n12712 = n1522 & n12695 ;
  assign n12649 = x[85] & n12633 ;
  assign n14370 = x[86] & n13533 ;
  assign n19135 = n12649 | n14370 ;
  assign n19136 = x[87] & n12631 ;
  assign n19137 = n19135 | n19136 ;
  assign n19138 = n12712 | n19137 ;
  assign n28744 = ~n19138 ;
  assign n19139 = x[11] & n28744 ;
  assign n19140 = n27892 & n19138 ;
  assign n19141 = n19139 | n19140 ;
  assign n28745 = ~n19141 ;
  assign n19142 = n19134 & n28745 ;
  assign n28746 = ~n19134 ;
  assign n19471 = n28746 & n19141 ;
  assign n19472 = n19142 | n19471 ;
  assign n19473 = n19470 & n19472 ;
  assign n20445 = n19470 | n19472 ;
  assign n28747 = ~n19473 ;
  assign n20446 = n28747 & n20445 ;
  assign n28748 = ~n20444 ;
  assign n20448 = n28748 & n20446 ;
  assign n28749 = ~n20446 ;
  assign n20449 = n20444 & n28749 ;
  assign n20450 = n20448 | n20449 ;
  assign n20460 = n20451 & n20458 ;
  assign n20813 = n20500 | n20812 ;
  assign n20814 = n20489 & n20813 ;
  assign n20815 = n20487 | n20814 ;
  assign n20817 = n20815 & n20816 ;
  assign n20818 = n20474 | n20817 ;
  assign n20819 = n20465 & n20818 ;
  assign n20820 = n20460 | n20819 ;
  assign n20821 = n20450 | n20820 ;
  assign n20822 = n20450 & n20820 ;
  assign n28750 = ~n20822 ;
  assign n21499 = n20821 & n28750 ;
  assign n18417 = n1685 & n18392 ;
  assign n18344 = x[91] & n18329 ;
  assign n18530 = x[92] & n18514 ;
  assign n21500 = n18344 | n18530 ;
  assign n21501 = x[93] & n18327 ;
  assign n21502 = n21500 | n21501 ;
  assign n21503 = n18417 | n21502 ;
  assign n28751 = ~n21503 ;
  assign n21504 = x[5] & n28751 ;
  assign n21505 = n27813 & n21503 ;
  assign n21506 = n21504 | n21505 ;
  assign n21507 = n21499 & n21506 ;
  assign n20447 = n20444 & n20446 ;
  assign n21128 = n20444 | n20446 ;
  assign n28752 = ~n20447 ;
  assign n21129 = n28752 & n21128 ;
  assign n28753 = ~n20820 ;
  assign n21130 = n28753 & n21129 ;
  assign n28754 = ~n21129 ;
  assign n22112 = n20820 & n28754 ;
  assign n22113 = n21130 | n22112 ;
  assign n22232 = n21506 | n22113 ;
  assign n28755 = ~n21507 ;
  assign n22943 = n28755 & n22232 ;
  assign n28756 = ~n22943 ;
  assign n22944 = n21935 & n28756 ;
  assign n22114 = n21506 & n22113 ;
  assign n22115 = n21516 & n21519 ;
  assign n22229 = n21533 | n22228 ;
  assign n22230 = n22116 & n22229 ;
  assign n22231 = n22115 | n22230 ;
  assign n22233 = n22231 & n22232 ;
  assign n22234 = n22114 | n22233 ;
  assign n28757 = ~n22234 ;
  assign n22945 = n22232 & n28757 ;
  assign n22946 = n22944 | n22945 ;
  assign n549 = n547 & n548 ;
  assign n550 = n27630 | n549 ;
  assign n25802 = x[95] & x[96] ;
  assign n551 = x[95] | x[96] ;
  assign n28758 = ~n25802 ;
  assign n1997 = n28758 & n551 ;
  assign n1998 = n550 & n1997 ;
  assign n1999 = n550 | n1997 ;
  assign n28759 = ~n1998 ;
  assign n2000 = n28759 & n1999 ;
  assign n19718 = n2000 & n19656 ;
  assign n19773 = x[94] & n19723 ;
  assign n19830 = x[95] & n19829 ;
  assign n22947 = n19773 | n19830 ;
  assign n22948 = x[96] & n19655 ;
  assign n22949 = n22947 | n22948 ;
  assign n22950 = n19718 | n22949 ;
  assign n28760 = ~n22950 ;
  assign n22951 = x[2] & n28760 ;
  assign n22952 = n27790 & n22950 ;
  assign n22953 = n22951 | n22952 ;
  assign n28761 = ~n22953 ;
  assign n22954 = n22946 & n28761 ;
  assign n28762 = ~n22946 ;
  assign n22955 = n28762 & n22953 ;
  assign n22956 = n22954 | n22955 ;
  assign n22957 = n22942 & n22956 ;
  assign n27669 = n22942 | n22956 ;
  assign n28763 = ~n22957 ;
  assign n161 = n28763 & n27669 ;
  assign n22958 = n22946 & n22953 ;
  assign n22959 = n22957 | n22958 ;
  assign n21936 = n21499 | n21506 ;
  assign n21937 = n21935 & n21936 ;
  assign n21938 = n21507 | n21937 ;
  assign n18412 = n2410 & n18392 ;
  assign n18391 = x[92] & n18329 ;
  assign n18532 = x[93] & n18514 ;
  assign n21490 = n18391 | n18532 ;
  assign n21491 = x[94] & n18327 ;
  assign n21492 = n21490 | n21491 ;
  assign n21493 = n18412 | n21492 ;
  assign n28764 = ~n21493 ;
  assign n21494 = x[5] & n28764 ;
  assign n21495 = n27813 & n21493 ;
  assign n21496 = n21494 | n21495 ;
  assign n15331 = n2046 & n15308 ;
  assign n15256 = x[89] & n15246 ;
  assign n17292 = x[90] & n16288 ;
  assign n20425 = n15256 | n17292 ;
  assign n20426 = x[91] & n15244 ;
  assign n20427 = n20425 | n20426 ;
  assign n20428 = n15331 | n20427 ;
  assign n28765 = ~n20428 ;
  assign n20429 = x[8] & n28765 ;
  assign n20430 = n27845 & n20428 ;
  assign n20431 = n20429 | n20430 ;
  assign n19143 = n19134 & n19141 ;
  assign n19474 = n19143 | n19473 ;
  assign n28766 = ~n16865 ;
  assign n16869 = n28766 & n16867 ;
  assign n28767 = ~n16867 ;
  assign n17759 = n16865 & n28767 ;
  assign n17760 = n16869 | n17759 ;
  assign n17802 = n17760 & n17800 ;
  assign n17803 = n16868 | n17802 ;
  assign n15962 = n15953 & n15960 ;
  assign n16447 = n15962 | n16446 ;
  assign n7219 = n1741 & n7162 ;
  assign n7108 = x[77] & n7100 ;
  assign n7723 = x[78] & n7647 ;
  assign n15940 = n7108 | n7723 ;
  assign n15941 = x[79] & n7098 ;
  assign n15942 = n15940 | n15941 ;
  assign n15943 = n7219 | n15942 ;
  assign n28768 = ~n15943 ;
  assign n15944 = x[20] & n28768 ;
  assign n15945 = n28114 & n15943 ;
  assign n15946 = n15944 | n15945 ;
  assign n15082 = n14932 | n14939 ;
  assign n15083 = n15081 & n15082 ;
  assign n15084 = n14940 | n15083 ;
  assign n14141 = n14041 | n14140 ;
  assign n5979 = n4632 & n5976 ;
  assign n4566 = x[68] & n4514 ;
  assign n4625 = x[69] & n4572 ;
  assign n13278 = n4566 | n4625 ;
  assign n13279 = x[70] & n4504 ;
  assign n13280 = n13278 | n13279 ;
  assign n13281 = n5979 | n13280 ;
  assign n28769 = ~n13281 ;
  assign n13282 = x[29] & n28769 ;
  assign n13283 = n28483 & n13281 ;
  assign n13284 = n13282 | n13283 ;
  assign n27737 = x[32] & x[33] ;
  assign n3902 = x[32] | x[33] ;
  assign n28770 = ~n27737 ;
  assign n3903 = n28770 & n3902 ;
  assign n11589 = x[64] & n3903 ;
  assign n12421 = n11589 & n28714 ;
  assign n28771 = ~n11589 ;
  assign n12422 = n28771 & n12420 ;
  assign n12423 = n12421 | n12422 ;
  assign n6504 = n779 & n6494 ;
  assign n672 = x[65] & n663 ;
  assign n753 = x[66] & n720 ;
  assign n12424 = n672 | n753 ;
  assign n12425 = x[67] & n652 ;
  assign n12426 = n12424 | n12425 ;
  assign n12427 = n6504 | n12426 ;
  assign n28772 = ~n12427 ;
  assign n12428 = x[32] & n28772 ;
  assign n12429 = n28658 & n12427 ;
  assign n12430 = n12428 | n12429 ;
  assign n28773 = ~n12430 ;
  assign n12431 = n12423 & n28773 ;
  assign n28774 = ~n12423 ;
  assign n13285 = n28774 & n12430 ;
  assign n13286 = n12431 | n13285 ;
  assign n28775 = ~n13284 ;
  assign n13287 = n28775 & n13286 ;
  assign n28776 = ~n13286 ;
  assign n13352 = n13284 & n28776 ;
  assign n13353 = n13287 | n13352 ;
  assign n28777 = ~n13353 ;
  assign n14018 = n13351 & n28777 ;
  assign n14019 = n28718 & n13353 ;
  assign n14020 = n14018 | n14019 ;
  assign n3735 = n452 & n3733 ;
  assign n338 = x[71] & n330 ;
  assign n421 = x[72] & n390 ;
  assign n14021 = n338 | n421 ;
  assign n14022 = x[73] & n322 ;
  assign n14023 = n14021 | n14022 ;
  assign n14024 = n3735 | n14023 ;
  assign n28778 = ~n14024 ;
  assign n14025 = x[26] & n28778 ;
  assign n14026 = n28342 & n14024 ;
  assign n14027 = n14025 | n14026 ;
  assign n14028 = n14020 | n14027 ;
  assign n14029 = n14020 & n14027 ;
  assign n28779 = ~n14029 ;
  assign n14142 = n14028 & n28779 ;
  assign n14143 = n14141 & n14142 ;
  assign n14921 = n14141 | n14142 ;
  assign n28780 = ~n14143 ;
  assign n14922 = n28780 & n14921 ;
  assign n5320 = n2750 & n5302 ;
  assign n5246 = x[74] & n5240 ;
  assign n6259 = x[75] & n6179 ;
  assign n14923 = n5246 | n6259 ;
  assign n14924 = x[76] & n5238 ;
  assign n14925 = n14923 | n14924 ;
  assign n14926 = n5320 | n14925 ;
  assign n28781 = ~n14926 ;
  assign n14927 = x[23] & n28781 ;
  assign n14928 = n28221 & n14926 ;
  assign n14929 = n14927 | n14928 ;
  assign n14930 = n14922 | n14929 ;
  assign n14931 = n14922 & n14929 ;
  assign n28782 = ~n14931 ;
  assign n15763 = n14930 & n28782 ;
  assign n28783 = ~n15084 ;
  assign n15765 = n28783 & n15763 ;
  assign n28784 = ~n15763 ;
  assign n15947 = n15084 & n28784 ;
  assign n15948 = n15765 | n15947 ;
  assign n28785 = ~n15946 ;
  assign n16147 = n28785 & n15948 ;
  assign n28786 = ~n15948 ;
  assign n16448 = n15946 & n28786 ;
  assign n16449 = n16147 | n16448 ;
  assign n16450 = n16447 | n16449 ;
  assign n16451 = n16447 & n16449 ;
  assign n28787 = ~n16451 ;
  assign n16849 = n16450 & n28787 ;
  assign n8713 = n1003 & n8706 ;
  assign n8657 = x[80] & n8645 ;
  assign n9890 = x[81] & n9278 ;
  assign n16850 = n8657 | n9890 ;
  assign n16851 = x[82] & n8643 ;
  assign n16852 = n16850 | n16851 ;
  assign n16853 = n8713 | n16852 ;
  assign n28788 = ~n16853 ;
  assign n16854 = x[17] & n28788 ;
  assign n16855 = n28039 & n16853 ;
  assign n16856 = n16854 | n16855 ;
  assign n16857 = n16849 | n16856 ;
  assign n16858 = n16849 & n16856 ;
  assign n28789 = ~n16858 ;
  assign n17804 = n16857 & n28789 ;
  assign n17805 = n17803 & n17804 ;
  assign n17878 = n17803 | n17804 ;
  assign n28790 = ~n17805 ;
  assign n17879 = n28790 & n17878 ;
  assign n10556 = n1239 & n10542 ;
  assign n10495 = x[83] & n10481 ;
  assign n11920 = x[84] & n11232 ;
  assign n17880 = n10495 | n11920 ;
  assign n17881 = x[85] & n10479 ;
  assign n17882 = n17880 | n17881 ;
  assign n17883 = n10556 | n17882 ;
  assign n28791 = ~n17883 ;
  assign n17884 = x[14] & n28791 ;
  assign n17885 = n27956 & n17883 ;
  assign n17886 = n17884 | n17885 ;
  assign n28792 = ~n17886 ;
  assign n17887 = n17879 & n28792 ;
  assign n28793 = ~n17879 ;
  assign n18181 = n28793 & n17886 ;
  assign n18182 = n17887 | n18181 ;
  assign n18183 = n18180 & n18182 ;
  assign n19049 = n18180 | n18182 ;
  assign n28794 = ~n18183 ;
  assign n19050 = n28794 & n19049 ;
  assign n12713 = n1720 & n12695 ;
  assign n12655 = x[86] & n12633 ;
  assign n14359 = x[87] & n13533 ;
  assign n19051 = n12655 | n14359 ;
  assign n19052 = x[88] & n12631 ;
  assign n19053 = n19051 | n19052 ;
  assign n19054 = n12713 | n19053 ;
  assign n28795 = ~n19054 ;
  assign n19055 = x[11] & n28795 ;
  assign n19056 = n27892 & n19054 ;
  assign n19057 = n19055 | n19056 ;
  assign n19058 = n19050 & n19057 ;
  assign n19475 = n19050 | n19057 ;
  assign n28796 = ~n19058 ;
  assign n20404 = n28796 & n19475 ;
  assign n28797 = ~n19474 ;
  assign n20406 = n28797 & n20404 ;
  assign n28798 = ~n20404 ;
  assign n20432 = n19474 & n28798 ;
  assign n20433 = n20406 | n20432 ;
  assign n28799 = ~n20431 ;
  assign n20435 = n28799 & n20433 ;
  assign n28800 = ~n20433 ;
  assign n21126 = n20431 & n28800 ;
  assign n21127 = n20435 | n21126 ;
  assign n21228 = n20464 | n21227 ;
  assign n21229 = n21129 & n21228 ;
  assign n21230 = n20447 | n21229 ;
  assign n21232 = n21127 | n21230 ;
  assign n21233 = n21127 & n21230 ;
  assign n28801 = ~n21233 ;
  assign n21939 = n21232 & n28801 ;
  assign n28802 = ~n21496 ;
  assign n21940 = n28802 & n21939 ;
  assign n28803 = ~n21939 ;
  assign n21941 = n21496 & n28803 ;
  assign n21942 = n21940 | n21941 ;
  assign n21943 = n21938 | n21942 ;
  assign n21944 = n21938 & n21942 ;
  assign n28804 = ~n21944 ;
  assign n22486 = n21943 & n28804 ;
  assign n552 = n550 & n551 ;
  assign n553 = n25802 | n552 ;
  assign n27628 = x[96] & x[97] ;
  assign n554 = x[96] | x[97] ;
  assign n28805 = ~n27628 ;
  assign n2435 = n28805 & n554 ;
  assign n2436 = n553 | n2435 ;
  assign n2437 = n553 & n2435 ;
  assign n28806 = ~n2437 ;
  assign n2438 = n2436 & n28806 ;
  assign n19695 = n2438 & n19656 ;
  assign n19741 = x[95] & n19723 ;
  assign n19865 = x[96] & n19829 ;
  assign n22487 = n19741 | n19865 ;
  assign n22488 = x[97] & n19655 ;
  assign n22489 = n22487 | n22488 ;
  assign n22490 = n19695 | n22489 ;
  assign n28807 = ~n22490 ;
  assign n22491 = x[2] & n28807 ;
  assign n22492 = n27790 & n22490 ;
  assign n22493 = n22491 | n22492 ;
  assign n22494 = n22486 | n22493 ;
  assign n22495 = n22486 & n22493 ;
  assign n28808 = ~n22495 ;
  assign n22960 = n22494 & n28808 ;
  assign n22961 = n22959 | n22960 ;
  assign n22962 = n22959 & n22960 ;
  assign n28809 = ~n22962 ;
  assign n162 = n22961 & n28809 ;
  assign n22963 = n22495 | n22962 ;
  assign n20434 = n20431 & n20433 ;
  assign n20436 = n20431 | n20433 ;
  assign n28810 = ~n20434 ;
  assign n20437 = n28810 & n20436 ;
  assign n28811 = ~n21230 ;
  assign n21231 = n20437 & n28811 ;
  assign n28812 = ~n20437 ;
  assign n21488 = n28812 & n21230 ;
  assign n21489 = n21231 | n21488 ;
  assign n21498 = n21489 & n21496 ;
  assign n21945 = n21498 | n21944 ;
  assign n19476 = n19474 & n19475 ;
  assign n19477 = n19058 | n19476 ;
  assign n8719 = n1057 & n8706 ;
  assign n8669 = x[81] & n8645 ;
  assign n9893 = x[82] & n9278 ;
  assign n16835 = n8669 | n9893 ;
  assign n16836 = x[83] & n8643 ;
  assign n16837 = n16835 | n16836 ;
  assign n16838 = n8719 | n16837 ;
  assign n28813 = ~n16838 ;
  assign n16839 = x[17] & n28813 ;
  assign n16840 = n28039 & n16838 ;
  assign n16841 = n16839 | n16840 ;
  assign n2723 = n452 & n2722 ;
  assign n340 = x[72] & n330 ;
  assign n444 = x[73] & n390 ;
  assign n14005 = n340 | n444 ;
  assign n14006 = x[74] & n322 ;
  assign n14007 = n14005 | n14006 ;
  assign n14008 = n2723 | n14007 ;
  assign n28814 = ~n14008 ;
  assign n14009 = x[26] & n28814 ;
  assign n14010 = n28342 & n14008 ;
  assign n14011 = n14009 | n14010 ;
  assign n13288 = n13284 & n13286 ;
  assign n13354 = n13351 & n13353 ;
  assign n13355 = n13288 | n13354 ;
  assign n4791 = n4632 & n4790 ;
  assign n4554 = x[69] & n4514 ;
  assign n4624 = x[70] & n4572 ;
  assign n13268 = n4554 | n4624 ;
  assign n13269 = x[71] & n4504 ;
  assign n13270 = n13268 | n13269 ;
  assign n13271 = n4791 | n13270 ;
  assign n28815 = ~n13271 ;
  assign n13272 = x[29] & n28815 ;
  assign n13273 = n28483 & n13271 ;
  assign n13274 = n13272 | n13273 ;
  assign n12432 = n12423 & n12430 ;
  assign n12433 = n11589 & n12420 ;
  assign n12434 = n12432 | n12433 ;
  assign n6410 = n779 & n6408 ;
  assign n678 = x[66] & n663 ;
  assign n772 = x[67] & n720 ;
  assign n12391 = n678 | n772 ;
  assign n12392 = x[68] & n652 ;
  assign n12393 = n12391 | n12392 ;
  assign n12394 = n6410 | n12393 ;
  assign n12395 = x[32] | n12394 ;
  assign n12396 = x[32] & n12394 ;
  assign n28816 = ~n12396 ;
  assign n12397 = n12395 & n28816 ;
  assign n11590 = x[35] & n28771 ;
  assign n27742 = x[34] & x[35] ;
  assign n3904 = x[34] | x[35] ;
  assign n28817 = ~n27742 ;
  assign n3905 = n28817 & n3904 ;
  assign n4041 = n3903 & n3905 ;
  assign n6444 = n4041 & n6437 ;
  assign n28818 = ~n3905 ;
  assign n3906 = n3903 & n28818 ;
  assign n11591 = x[65] & n3906 ;
  assign n27747 = x[33] & x[34] ;
  assign n3907 = x[33] | x[34] ;
  assign n28819 = ~n27747 ;
  assign n3908 = n28819 & n3907 ;
  assign n28820 = ~n3903 ;
  assign n3975 = n28820 & n3908 ;
  assign n11592 = x[64] & n3975 ;
  assign n11593 = n11591 | n11592 ;
  assign n11594 = n6444 | n11593 ;
  assign n28821 = ~n11594 ;
  assign n11595 = x[35] & n28821 ;
  assign n28822 = ~x[35] ;
  assign n11596 = n28822 & n11594 ;
  assign n11597 = n11595 | n11596 ;
  assign n28823 = ~n11597 ;
  assign n11598 = n11590 & n28823 ;
  assign n28824 = ~n11590 ;
  assign n12398 = n28824 & n11597 ;
  assign n12399 = n11598 | n12398 ;
  assign n12400 = n12397 & n12399 ;
  assign n12435 = n12397 | n12399 ;
  assign n28825 = ~n12400 ;
  assign n12436 = n28825 & n12435 ;
  assign n28826 = ~n12434 ;
  assign n12437 = n28826 & n12436 ;
  assign n28827 = ~n12436 ;
  assign n13275 = n12434 & n28827 ;
  assign n13276 = n12437 | n13275 ;
  assign n13277 = n13274 | n13276 ;
  assign n13356 = n13274 & n13276 ;
  assign n28828 = ~n13356 ;
  assign n13357 = n13277 & n28828 ;
  assign n13358 = n13355 & n13357 ;
  assign n14012 = n13355 | n13357 ;
  assign n28829 = ~n13358 ;
  assign n14013 = n28829 & n14012 ;
  assign n28830 = ~n14011 ;
  assign n14014 = n28830 & n14013 ;
  assign n28831 = ~n14013 ;
  assign n14016 = n14011 & n28831 ;
  assign n14017 = n14014 | n14016 ;
  assign n14144 = n14029 | n14143 ;
  assign n14145 = n14017 | n14144 ;
  assign n14147 = n14017 & n14144 ;
  assign n28832 = ~n14147 ;
  assign n14912 = n14145 & n28832 ;
  assign n5303 = n1775 & n5302 ;
  assign n5289 = x[75] & n5240 ;
  assign n6227 = x[76] & n6179 ;
  assign n14913 = n5289 | n6227 ;
  assign n14914 = x[77] & n5238 ;
  assign n14915 = n14913 | n14914 ;
  assign n14916 = n5303 | n14915 ;
  assign n28833 = ~n14916 ;
  assign n14917 = x[23] & n28833 ;
  assign n14918 = n28221 & n14916 ;
  assign n14919 = n14917 | n14918 ;
  assign n15087 = n14912 | n14919 ;
  assign n14920 = n14912 & n14919 ;
  assign n15085 = n14930 & n15084 ;
  assign n15086 = n14931 | n15085 ;
  assign n15088 = n15086 & n15087 ;
  assign n15089 = n14920 | n15088 ;
  assign n28834 = ~n15089 ;
  assign n15090 = n15087 & n28834 ;
  assign n28835 = ~n14144 ;
  assign n14146 = n14017 & n28835 ;
  assign n28836 = ~n14017 ;
  assign n15739 = n28836 & n14144 ;
  assign n15740 = n14146 | n15739 ;
  assign n15741 = n14919 & n15740 ;
  assign n28837 = ~n15741 ;
  assign n15742 = n15087 & n28837 ;
  assign n15764 = n15762 & n15763 ;
  assign n15766 = n14931 | n15764 ;
  assign n28838 = ~n15742 ;
  assign n15928 = n28838 & n15766 ;
  assign n15929 = n15090 | n15928 ;
  assign n7171 = n1270 & n7162 ;
  assign n7109 = x[78] & n7100 ;
  assign n7682 = x[79] & n7647 ;
  assign n15930 = n7109 | n7682 ;
  assign n15931 = x[80] & n7098 ;
  assign n15932 = n15930 | n15931 ;
  assign n15933 = n7171 | n15932 ;
  assign n28839 = ~n15933 ;
  assign n15934 = x[20] & n28839 ;
  assign n15935 = n28114 & n15933 ;
  assign n15936 = n15934 | n15935 ;
  assign n15937 = n15929 | n15936 ;
  assign n15938 = n15929 & n15936 ;
  assign n28840 = ~n15938 ;
  assign n15939 = n15937 & n28840 ;
  assign n15949 = n15946 & n15948 ;
  assign n15972 = n15963 & n15970 ;
  assign n16140 = n16138 & n16139 ;
  assign n16141 = n15987 | n16140 ;
  assign n16142 = n15977 & n16141 ;
  assign n16143 = n15972 | n16142 ;
  assign n16144 = n15953 | n15960 ;
  assign n16145 = n16143 & n16144 ;
  assign n16146 = n15962 | n16145 ;
  assign n16148 = n15946 | n15948 ;
  assign n28841 = ~n15949 ;
  assign n16149 = n28841 & n16148 ;
  assign n16150 = n16146 & n16149 ;
  assign n16151 = n15949 | n16150 ;
  assign n28842 = ~n16151 ;
  assign n16420 = n15939 & n28842 ;
  assign n28843 = ~n15939 ;
  assign n16844 = n28843 & n16151 ;
  assign n16845 = n16420 | n16844 ;
  assign n16846 = n16841 | n16845 ;
  assign n16847 = n16841 & n16845 ;
  assign n28844 = ~n16847 ;
  assign n16848 = n16846 & n28844 ;
  assign n17806 = n16858 | n17805 ;
  assign n28845 = ~n17806 ;
  assign n17807 = n16848 & n28845 ;
  assign n28846 = ~n16848 ;
  assign n17866 = n28846 & n17806 ;
  assign n17867 = n17807 | n17866 ;
  assign n10560 = n1213 & n10542 ;
  assign n10539 = x[84] & n10481 ;
  assign n11917 = x[85] & n11232 ;
  assign n17868 = n10539 | n11917 ;
  assign n17869 = x[86] & n10479 ;
  assign n17870 = n17868 | n17869 ;
  assign n17871 = n10560 | n17870 ;
  assign n28847 = ~n17871 ;
  assign n17872 = x[14] & n28847 ;
  assign n17873 = n27956 & n17871 ;
  assign n17874 = n17872 | n17873 ;
  assign n17875 = n17867 | n17874 ;
  assign n17876 = n17867 & n17874 ;
  assign n28848 = ~n17876 ;
  assign n17877 = n17875 & n28848 ;
  assign n17888 = n17879 & n17886 ;
  assign n18184 = n17888 | n18183 ;
  assign n28849 = ~n18184 ;
  assign n18185 = n17877 & n28849 ;
  assign n28850 = ~n17877 ;
  assign n19039 = n28850 & n18184 ;
  assign n19040 = n18185 | n19039 ;
  assign n12714 = n1453 & n12695 ;
  assign n12651 = x[87] & n12633 ;
  assign n14373 = x[88] & n13533 ;
  assign n19041 = n12651 | n14373 ;
  assign n19042 = x[89] & n12631 ;
  assign n19043 = n19041 | n19042 ;
  assign n19044 = n12714 | n19043 ;
  assign n28851 = ~n19044 ;
  assign n19045 = x[11] & n28851 ;
  assign n19046 = n27892 & n19044 ;
  assign n19047 = n19045 | n19046 ;
  assign n19048 = n19040 & n19047 ;
  assign n19478 = n19040 | n19047 ;
  assign n28852 = ~n19048 ;
  assign n20410 = n28852 & n19478 ;
  assign n28853 = ~n20410 ;
  assign n20411 = n19477 & n28853 ;
  assign n20319 = n19152 & n19156 ;
  assign n20398 = n19464 | n20397 ;
  assign n20399 = n20320 & n20398 ;
  assign n20400 = n20319 | n20399 ;
  assign n20401 = n19134 | n19141 ;
  assign n20402 = n20400 & n20401 ;
  assign n20403 = n19143 | n20402 ;
  assign n20405 = n20403 & n20404 ;
  assign n20407 = n19058 | n20405 ;
  assign n20408 = n19478 & n20407 ;
  assign n20409 = n19048 | n20408 ;
  assign n28854 = ~n20409 ;
  assign n20412 = n19478 & n28854 ;
  assign n20413 = n20411 | n20412 ;
  assign n15334 = n1841 & n15308 ;
  assign n15286 = x[90] & n15246 ;
  assign n17296 = x[91] & n16288 ;
  assign n20414 = n15286 | n17296 ;
  assign n20415 = x[92] & n15244 ;
  assign n20416 = n20414 | n20415 ;
  assign n20417 = n15334 | n20416 ;
  assign n28855 = ~n20417 ;
  assign n20418 = x[8] & n28855 ;
  assign n20419 = n27845 & n20417 ;
  assign n20420 = n20418 | n20419 ;
  assign n28856 = ~n20420 ;
  assign n20421 = n20413 & n28856 ;
  assign n28857 = ~n20413 ;
  assign n20423 = n28857 & n20420 ;
  assign n20424 = n20421 | n20423 ;
  assign n20823 = n20447 | n20822 ;
  assign n20824 = n20437 & n20823 ;
  assign n20825 = n20434 | n20824 ;
  assign n20826 = n20424 | n20825 ;
  assign n20827 = n20424 & n20825 ;
  assign n28858 = ~n20827 ;
  assign n21479 = n20826 & n28858 ;
  assign n18413 = n2152 & n18392 ;
  assign n18346 = x[93] & n18329 ;
  assign n18534 = x[94] & n18514 ;
  assign n21480 = n18346 | n18534 ;
  assign n21481 = x[95] & n18327 ;
  assign n21482 = n21480 | n21481 ;
  assign n21483 = n18413 | n21482 ;
  assign n28859 = ~n21483 ;
  assign n21484 = x[5] & n28859 ;
  assign n21485 = n27813 & n21483 ;
  assign n21486 = n21484 | n21485 ;
  assign n21487 = n21479 & n21486 ;
  assign n28860 = ~n20825 ;
  assign n21125 = n20424 & n28860 ;
  assign n28861 = ~n20424 ;
  assign n22108 = n28861 & n20825 ;
  assign n22109 = n21125 | n22108 ;
  assign n22238 = n21486 | n22109 ;
  assign n28862 = ~n21487 ;
  assign n22964 = n28862 & n22238 ;
  assign n28863 = ~n22964 ;
  assign n22965 = n21945 & n28863 ;
  assign n22110 = n21486 & n22109 ;
  assign n22111 = n21496 & n21939 ;
  assign n21497 = n21489 | n21496 ;
  assign n28864 = ~n21498 ;
  assign n22235 = n21497 & n28864 ;
  assign n22236 = n22234 & n22235 ;
  assign n22237 = n22111 | n22236 ;
  assign n22239 = n22237 & n22238 ;
  assign n22240 = n22110 | n22239 ;
  assign n28865 = ~n22240 ;
  assign n22966 = n22238 & n28865 ;
  assign n22967 = n22965 | n22966 ;
  assign n555 = n553 & n554 ;
  assign n556 = n27628 | n555 ;
  assign n25668 = x[97] & x[98] ;
  assign n557 = x[97] | x[98] ;
  assign n28866 = ~n25668 ;
  assign n2838 = n28866 & n557 ;
  assign n2839 = n556 & n2838 ;
  assign n2840 = n556 | n2838 ;
  assign n28867 = ~n2839 ;
  assign n2841 = n28867 & n2840 ;
  assign n19719 = n2841 & n19656 ;
  assign n19785 = x[96] & n19723 ;
  assign n19890 = x[97] & n19829 ;
  assign n22968 = n19785 | n19890 ;
  assign n22969 = x[98] & n19655 ;
  assign n22970 = n22968 | n22969 ;
  assign n22971 = n19719 | n22970 ;
  assign n28868 = ~n22971 ;
  assign n22972 = x[2] & n28868 ;
  assign n22973 = n27790 & n22971 ;
  assign n22974 = n22972 | n22973 ;
  assign n28869 = ~n22974 ;
  assign n22975 = n22967 & n28869 ;
  assign n28870 = ~n22967 ;
  assign n22976 = n28870 & n22974 ;
  assign n22977 = n22975 | n22976 ;
  assign n22978 = n22963 & n22977 ;
  assign n27672 = n22963 | n22977 ;
  assign n28871 = ~n22978 ;
  assign n163 = n28871 & n27672 ;
  assign n22979 = n22967 & n22974 ;
  assign n22980 = n22978 | n22979 ;
  assign n18414 = n2000 & n18392 ;
  assign n18347 = x[94] & n18329 ;
  assign n18535 = x[95] & n18514 ;
  assign n21471 = n18347 | n18535 ;
  assign n21472 = x[96] & n18327 ;
  assign n21473 = n21471 | n21472 ;
  assign n21474 = n18414 | n21473 ;
  assign n28872 = ~n21474 ;
  assign n21475 = x[5] & n28872 ;
  assign n21476 = n27813 & n21474 ;
  assign n21477 = n21475 | n21476 ;
  assign n15335 = n1685 & n15308 ;
  assign n15292 = x[91] & n15246 ;
  assign n17306 = x[92] & n16288 ;
  assign n20306 = n15292 | n17306 ;
  assign n20307 = x[93] & n15244 ;
  assign n20308 = n20306 | n20307 ;
  assign n20309 = n15335 | n20308 ;
  assign n28873 = ~n20309 ;
  assign n20310 = x[8] & n28873 ;
  assign n20311 = n27845 & n20309 ;
  assign n20312 = n20310 | n20311 ;
  assign n19479 = n19477 & n19478 ;
  assign n19480 = n19048 | n19479 ;
  assign n12715 = n1482 & n12695 ;
  assign n12642 = x[88] & n12633 ;
  assign n14403 = x[89] & n13533 ;
  assign n19029 = n12642 | n14403 ;
  assign n19030 = x[90] & n12631 ;
  assign n19031 = n19029 | n19030 ;
  assign n19032 = n12715 | n19031 ;
  assign n19033 = x[11] | n19032 ;
  assign n19034 = x[11] & n19032 ;
  assign n28874 = ~n19034 ;
  assign n19035 = n19033 & n28874 ;
  assign n18186 = n17877 & n18184 ;
  assign n18187 = n17876 | n18186 ;
  assign n16152 = n15939 | n16151 ;
  assign n16153 = n15939 & n16151 ;
  assign n28875 = ~n16153 ;
  assign n16834 = n16152 & n28875 ;
  assign n28876 = ~n16841 ;
  assign n16842 = n16834 & n28876 ;
  assign n28877 = ~n16834 ;
  assign n17757 = n28877 & n16841 ;
  assign n17758 = n16842 | n17757 ;
  assign n17808 = n17758 & n17806 ;
  assign n17809 = n16847 | n17808 ;
  assign n7180 = n1029 & n7162 ;
  assign n7110 = x[79] & n7100 ;
  assign n7706 = x[80] & n7647 ;
  assign n15915 = n7110 | n7706 ;
  assign n15916 = x[81] & n7098 ;
  assign n15917 = n15915 | n15916 ;
  assign n15918 = n7180 | n15917 ;
  assign n28878 = ~n15918 ;
  assign n15919 = x[20] & n28878 ;
  assign n15920 = n28114 & n15918 ;
  assign n15921 = n15919 | n15920 ;
  assign n15767 = n14919 | n15740 ;
  assign n15768 = n15766 & n15767 ;
  assign n15769 = n15741 | n15768 ;
  assign n14015 = n14011 & n14013 ;
  assign n14148 = n14015 | n14147 ;
  assign n3292 = n452 & n3289 ;
  assign n352 = x[73] & n330 ;
  assign n402 = x[74] & n390 ;
  assign n13995 = n352 | n402 ;
  assign n13996 = x[75] & n322 ;
  assign n13997 = n13995 | n13996 ;
  assign n13998 = n3292 | n13997 ;
  assign n28879 = ~n13998 ;
  assign n13999 = x[26] & n28879 ;
  assign n14000 = n28342 & n13998 ;
  assign n14001 = n13999 | n14000 ;
  assign n13359 = n13356 | n13358 ;
  assign n12438 = n12434 & n12436 ;
  assign n12439 = n12400 | n12438 ;
  assign n11599 = n11590 & n11597 ;
  assign n6468 = n4041 & n6466 ;
  assign n3909 = n28820 & n3905 ;
  assign n28880 = ~n3908 ;
  assign n3910 = n28880 & n3909 ;
  assign n3944 = x[64] & n3910 ;
  assign n3979 = x[65] & n3975 ;
  assign n11600 = n3944 | n3979 ;
  assign n11601 = x[66] & n3906 ;
  assign n11602 = n11600 | n11601 ;
  assign n11603 = n6468 | n11602 ;
  assign n28881 = ~n11603 ;
  assign n11604 = x[35] & n28881 ;
  assign n11605 = n28822 & n11603 ;
  assign n11606 = n11604 | n11605 ;
  assign n11607 = n11599 | n11606 ;
  assign n11608 = n11599 & n11606 ;
  assign n28882 = ~n11608 ;
  assign n12382 = n11607 & n28882 ;
  assign n6383 = n779 & n6379 ;
  assign n717 = x[67] & n663 ;
  assign n770 = x[68] & n720 ;
  assign n12383 = n717 | n770 ;
  assign n12384 = x[69] & n652 ;
  assign n12385 = n12383 | n12384 ;
  assign n12386 = n6383 | n12385 ;
  assign n28883 = ~n12386 ;
  assign n12387 = x[32] & n28883 ;
  assign n12388 = n28658 & n12386 ;
  assign n12389 = n12387 | n12388 ;
  assign n12390 = n12382 & n12389 ;
  assign n12440 = n12382 | n12389 ;
  assign n28884 = ~n12390 ;
  assign n13255 = n28884 & n12440 ;
  assign n28885 = ~n13255 ;
  assign n13256 = n12439 & n28885 ;
  assign n12441 = n12439 & n12440 ;
  assign n12442 = n12390 | n12441 ;
  assign n28886 = ~n12442 ;
  assign n13257 = n12440 & n28886 ;
  assign n13258 = n13256 | n13257 ;
  assign n4633 = n3701 & n4632 ;
  assign n4565 = x[70] & n4514 ;
  assign n4614 = x[71] & n4572 ;
  assign n13259 = n4565 | n4614 ;
  assign n13260 = x[72] & n4504 ;
  assign n13261 = n13259 | n13260 ;
  assign n13262 = n4633 | n13261 ;
  assign n28887 = ~n13262 ;
  assign n13263 = x[29] & n28887 ;
  assign n13264 = n28483 & n13262 ;
  assign n13265 = n13263 | n13264 ;
  assign n28888 = ~n13265 ;
  assign n13266 = n13258 & n28888 ;
  assign n28889 = ~n13258 ;
  assign n13360 = n28889 & n13265 ;
  assign n13361 = n13266 | n13360 ;
  assign n28890 = ~n13361 ;
  assign n13362 = n13359 & n28890 ;
  assign n28891 = ~n13359 ;
  assign n14002 = n28891 & n13361 ;
  assign n14003 = n13362 | n14002 ;
  assign n28892 = ~n14001 ;
  assign n14149 = n28892 & n14003 ;
  assign n28893 = ~n14003 ;
  assign n14712 = n14001 & n28893 ;
  assign n14713 = n14149 | n14712 ;
  assign n28894 = ~n14713 ;
  assign n14714 = n14148 & n28894 ;
  assign n28895 = ~n14148 ;
  assign n14901 = n28895 & n14713 ;
  assign n14902 = n14714 | n14901 ;
  assign n5323 = n2084 & n5302 ;
  assign n5247 = x[76] & n5240 ;
  assign n6245 = x[77] & n6179 ;
  assign n14903 = n5247 | n6245 ;
  assign n14904 = x[78] & n5238 ;
  assign n14905 = n14903 | n14904 ;
  assign n14906 = n5323 | n14905 ;
  assign n28896 = ~n14906 ;
  assign n14907 = x[23] & n28896 ;
  assign n14908 = n28221 & n14906 ;
  assign n14909 = n14907 | n14908 ;
  assign n14910 = n14902 | n14909 ;
  assign n14911 = n14902 & n14909 ;
  assign n28897 = ~n14911 ;
  assign n15770 = n14910 & n28897 ;
  assign n15771 = n15769 & n15770 ;
  assign n15922 = n15769 | n15770 ;
  assign n28898 = ~n15771 ;
  assign n15923 = n28898 & n15922 ;
  assign n15924 = n15921 & n15923 ;
  assign n15926 = n15921 | n15923 ;
  assign n28899 = ~n15924 ;
  assign n15927 = n28899 & n15926 ;
  assign n16452 = n15949 | n16451 ;
  assign n16453 = n15939 & n16452 ;
  assign n16454 = n15938 | n16453 ;
  assign n28900 = ~n16454 ;
  assign n16455 = n15927 & n28900 ;
  assign n28901 = ~n15927 ;
  assign n16824 = n28901 & n16454 ;
  assign n16825 = n16455 | n16824 ;
  assign n8709 = n1293 & n8706 ;
  assign n8654 = x[82] & n8645 ;
  assign n9891 = x[83] & n9278 ;
  assign n16826 = n8654 | n9891 ;
  assign n16827 = x[84] & n8643 ;
  assign n16828 = n16826 | n16827 ;
  assign n16829 = n8709 | n16828 ;
  assign n28902 = ~n16829 ;
  assign n16830 = x[17] & n28902 ;
  assign n16831 = n28039 & n16829 ;
  assign n16832 = n16830 | n16831 ;
  assign n17111 = n16825 | n16832 ;
  assign n28903 = ~n15921 ;
  assign n15925 = n28903 & n15923 ;
  assign n28904 = ~n15923 ;
  assign n16418 = n15921 & n28904 ;
  assign n16419 = n15925 | n16418 ;
  assign n16456 = n16419 | n16454 ;
  assign n16457 = n16419 & n16454 ;
  assign n28905 = ~n16457 ;
  assign n17755 = n16456 & n28905 ;
  assign n17756 = n16832 & n17755 ;
  assign n28906 = ~n17756 ;
  assign n17853 = n17111 & n28906 ;
  assign n28907 = ~n17853 ;
  assign n17854 = n17809 & n28907 ;
  assign n16833 = n16825 & n16832 ;
  assign n16843 = n16834 & n16841 ;
  assign n28908 = ~n16878 ;
  assign n16883 = n28908 & n16882 ;
  assign n28909 = ~n16882 ;
  assign n16885 = n16878 & n28909 ;
  assign n16886 = n16883 | n16885 ;
  assign n17103 = n16886 & n17102 ;
  assign n17104 = n16881 | n17103 ;
  assign n17105 = n16871 & n17104 ;
  assign n17106 = n16868 | n17105 ;
  assign n17107 = n16857 & n17106 ;
  assign n17108 = n16858 | n17107 ;
  assign n17109 = n16848 & n17108 ;
  assign n17110 = n16843 | n17109 ;
  assign n17112 = n17110 & n17111 ;
  assign n17113 = n16833 | n17112 ;
  assign n28910 = ~n17113 ;
  assign n17855 = n17111 & n28910 ;
  assign n17856 = n17854 | n17855 ;
  assign n10592 = n1522 & n10542 ;
  assign n10499 = x[85] & n10481 ;
  assign n11916 = x[86] & n11232 ;
  assign n17857 = n10499 | n11916 ;
  assign n17858 = x[87] & n10479 ;
  assign n17859 = n17857 | n17858 ;
  assign n17860 = n10592 | n17859 ;
  assign n28911 = ~n17860 ;
  assign n17861 = x[14] & n28911 ;
  assign n17862 = n27956 & n17860 ;
  assign n17863 = n17861 | n17862 ;
  assign n28912 = ~n17863 ;
  assign n17864 = n17856 & n28912 ;
  assign n28913 = ~n17856 ;
  assign n18188 = n28913 & n17863 ;
  assign n18189 = n17864 | n18188 ;
  assign n18190 = n18187 & n18189 ;
  assign n19036 = n18187 | n18189 ;
  assign n28914 = ~n18190 ;
  assign n19037 = n28914 & n19036 ;
  assign n19038 = n19035 & n19037 ;
  assign n19481 = n19035 | n19037 ;
  assign n28915 = ~n19038 ;
  assign n19482 = n28915 & n19481 ;
  assign n28916 = ~n19480 ;
  assign n19483 = n28916 & n19482 ;
  assign n28917 = ~n19482 ;
  assign n20313 = n19480 & n28917 ;
  assign n20314 = n19483 | n20313 ;
  assign n28918 = ~n20312 ;
  assign n20316 = n28918 & n20314 ;
  assign n28919 = ~n20314 ;
  assign n21123 = n20312 & n28919 ;
  assign n21124 = n20316 | n21123 ;
  assign n20422 = n20413 & n20420 ;
  assign n21234 = n20434 | n21233 ;
  assign n21235 = n20424 & n21234 ;
  assign n21236 = n20422 | n21235 ;
  assign n21238 = n21124 | n21236 ;
  assign n21239 = n21124 & n21236 ;
  assign n28920 = ~n21239 ;
  assign n22106 = n21238 & n28920 ;
  assign n22241 = n21477 | n22106 ;
  assign n22107 = n21477 & n22106 ;
  assign n22242 = n22240 & n22241 ;
  assign n22244 = n22107 | n22242 ;
  assign n28921 = ~n22244 ;
  assign n22245 = n22241 & n28921 ;
  assign n21946 = n21479 | n21486 ;
  assign n21947 = n21945 & n21946 ;
  assign n21948 = n21487 | n21947 ;
  assign n20315 = n20312 & n20314 ;
  assign n20317 = n20312 | n20314 ;
  assign n28922 = ~n20315 ;
  assign n20318 = n28922 & n20317 ;
  assign n28923 = ~n21236 ;
  assign n21237 = n20318 & n28923 ;
  assign n28924 = ~n20318 ;
  assign n21469 = n28924 & n21236 ;
  assign n21470 = n21237 | n21469 ;
  assign n21478 = n21470 & n21477 ;
  assign n28925 = ~n21478 ;
  assign n22243 = n28925 & n22241 ;
  assign n28926 = ~n22243 ;
  assign n22981 = n21948 & n28926 ;
  assign n22982 = n22245 | n22981 ;
  assign n558 = n556 & n557 ;
  assign n559 = n25668 | n558 ;
  assign n27627 = x[98] & x[99] ;
  assign n560 = x[98] | x[99] ;
  assign n28927 = ~n27627 ;
  assign n2310 = n28927 & n560 ;
  assign n2311 = n559 | n2310 ;
  assign n2312 = n559 & n2310 ;
  assign n28928 = ~n2312 ;
  assign n2313 = n2311 & n28928 ;
  assign n19720 = n2313 & n19656 ;
  assign n19786 = x[97] & n19723 ;
  assign n19838 = x[98] & n19829 ;
  assign n22983 = n19786 | n19838 ;
  assign n22984 = x[99] & n19655 ;
  assign n22985 = n22983 | n22984 ;
  assign n22986 = n19720 | n22985 ;
  assign n28929 = ~n22986 ;
  assign n22987 = x[2] & n28929 ;
  assign n22988 = n27790 & n22986 ;
  assign n22989 = n22987 | n22988 ;
  assign n22990 = n22982 | n22989 ;
  assign n22991 = n22982 & n22989 ;
  assign n28930 = ~n22991 ;
  assign n22992 = n22990 & n28930 ;
  assign n22993 = n22980 | n22992 ;
  assign n22994 = n22980 & n22992 ;
  assign n28931 = ~n22994 ;
  assign n164 = n22993 & n28931 ;
  assign n21949 = n21470 | n21477 ;
  assign n21950 = n21948 & n21949 ;
  assign n21951 = n21478 | n21950 ;
  assign n18415 = n2438 & n18392 ;
  assign n18351 = x[95] & n18329 ;
  assign n18547 = x[96] & n18514 ;
  assign n21459 = n18351 | n18547 ;
  assign n21460 = x[97] & n18327 ;
  assign n21461 = n21459 | n21460 ;
  assign n21462 = n18415 | n21461 ;
  assign n28932 = ~n21462 ;
  assign n21463 = x[5] & n28932 ;
  assign n21464 = n27813 & n21462 ;
  assign n21465 = n21463 | n21464 ;
  assign n21240 = n20315 | n21239 ;
  assign n19484 = n19480 & n19482 ;
  assign n19485 = n19038 | n19484 ;
  assign n12723 = n2046 & n12695 ;
  assign n12668 = x[89] & n12633 ;
  assign n14354 = x[90] & n13533 ;
  assign n19019 = n12668 | n14354 ;
  assign n19020 = x[91] & n12631 ;
  assign n19021 = n19019 | n19020 ;
  assign n19022 = n12723 | n19021 ;
  assign n28933 = ~n19022 ;
  assign n19023 = x[11] & n28933 ;
  assign n19024 = n27892 & n19022 ;
  assign n19025 = n19023 | n19024 ;
  assign n17865 = n17856 & n17863 ;
  assign n18191 = n17865 | n18190 ;
  assign n17810 = n16832 | n17755 ;
  assign n17811 = n17809 & n17810 ;
  assign n17812 = n17756 | n17811 ;
  assign n16458 = n15924 | n16457 ;
  assign n15772 = n14911 | n15771 ;
  assign n5304 = n1741 & n5302 ;
  assign n5293 = x[77] & n5240 ;
  assign n6265 = x[78] & n6179 ;
  assign n14891 = n5293 | n6265 ;
  assign n14892 = x[79] & n5238 ;
  assign n14893 = n14891 | n14892 ;
  assign n14894 = n5304 | n14893 ;
  assign n28934 = ~n14894 ;
  assign n14895 = x[23] & n28934 ;
  assign n14896 = n28221 & n14894 ;
  assign n14897 = n14895 | n14896 ;
  assign n2751 = n452 & n2750 ;
  assign n368 = x[74] & n330 ;
  assign n443 = x[75] & n390 ;
  assign n13981 = n368 | n443 ;
  assign n13982 = x[76] & n322 ;
  assign n13983 = n13981 | n13982 ;
  assign n13984 = n2751 | n13983 ;
  assign n28935 = ~n13984 ;
  assign n13985 = x[26] & n28935 ;
  assign n13986 = n28342 & n13984 ;
  assign n13987 = n13985 | n13986 ;
  assign n13267 = n13258 & n13265 ;
  assign n13363 = n13359 & n13361 ;
  assign n13364 = n13267 | n13363 ;
  assign n5986 = n779 & n5976 ;
  assign n715 = x[68] & n663 ;
  assign n751 = x[69] & n720 ;
  assign n12371 = n715 | n751 ;
  assign n12372 = x[70] & n652 ;
  assign n12373 = n12371 | n12372 ;
  assign n12374 = n5986 | n12373 ;
  assign n28936 = ~n12374 ;
  assign n12375 = x[32] & n28936 ;
  assign n12376 = n28658 & n12374 ;
  assign n12377 = n12375 | n12376 ;
  assign n27728 = x[35] & x[36] ;
  assign n3435 = x[35] | x[36] ;
  assign n28937 = ~n27728 ;
  assign n3436 = n28937 & n3435 ;
  assign n10992 = x[64] & n3436 ;
  assign n11609 = n10992 & n28882 ;
  assign n28938 = ~n10992 ;
  assign n11610 = n28938 & n11608 ;
  assign n11611 = n11609 | n11610 ;
  assign n6496 = n4041 & n6494 ;
  assign n3918 = x[65] & n3910 ;
  assign n3978 = x[66] & n3975 ;
  assign n11612 = n3918 | n3978 ;
  assign n11613 = x[67] & n3906 ;
  assign n11614 = n11612 | n11613 ;
  assign n11615 = n6496 | n11614 ;
  assign n28939 = ~n11615 ;
  assign n11616 = x[35] & n28939 ;
  assign n11617 = n28822 & n11615 ;
  assign n11618 = n11616 | n11617 ;
  assign n28940 = ~n11618 ;
  assign n11619 = n11611 & n28940 ;
  assign n28941 = ~n11611 ;
  assign n12378 = n28941 & n11618 ;
  assign n12379 = n11619 | n12378 ;
  assign n28942 = ~n12377 ;
  assign n12380 = n28942 & n12379 ;
  assign n28943 = ~n12379 ;
  assign n12443 = n12377 & n28943 ;
  assign n12444 = n12380 | n12443 ;
  assign n28944 = ~n12444 ;
  assign n13243 = n12442 & n28944 ;
  assign n13244 = n28886 & n12444 ;
  assign n13245 = n13243 | n13244 ;
  assign n4645 = n3733 & n4632 ;
  assign n4564 = x[71] & n4514 ;
  assign n4623 = x[72] & n4572 ;
  assign n13246 = n4564 | n4623 ;
  assign n13247 = x[73] & n4504 ;
  assign n13248 = n13246 | n13247 ;
  assign n13249 = n4645 | n13248 ;
  assign n28945 = ~n13249 ;
  assign n13250 = x[29] & n28945 ;
  assign n13251 = n28483 & n13249 ;
  assign n13252 = n13250 | n13251 ;
  assign n13253 = n13245 | n13252 ;
  assign n13254 = n13245 & n13252 ;
  assign n28946 = ~n13254 ;
  assign n13365 = n13253 & n28946 ;
  assign n13366 = n13364 & n13365 ;
  assign n13990 = n13364 | n13365 ;
  assign n28947 = ~n13366 ;
  assign n13991 = n28947 & n13990 ;
  assign n28948 = ~n13987 ;
  assign n13992 = n28948 & n13991 ;
  assign n28949 = ~n13991 ;
  assign n13993 = n13987 & n28949 ;
  assign n13994 = n13992 | n13993 ;
  assign n14004 = n14001 & n14003 ;
  assign n14150 = n14001 | n14003 ;
  assign n28950 = ~n14004 ;
  assign n14151 = n28950 & n14150 ;
  assign n14152 = n14148 & n14151 ;
  assign n14153 = n14004 | n14152 ;
  assign n14154 = n13994 | n14153 ;
  assign n14155 = n13994 & n14153 ;
  assign n28951 = ~n14155 ;
  assign n15093 = n14154 & n28951 ;
  assign n28952 = ~n14897 ;
  assign n15095 = n28952 & n15093 ;
  assign n28953 = ~n15093 ;
  assign n15773 = n14897 & n28953 ;
  assign n15774 = n15095 | n15773 ;
  assign n15775 = n15772 | n15774 ;
  assign n15776 = n15772 & n15774 ;
  assign n28954 = ~n15776 ;
  assign n15906 = n15775 & n28954 ;
  assign n7194 = n1003 & n7162 ;
  assign n7122 = x[80] & n7100 ;
  assign n7683 = x[81] & n7647 ;
  assign n15907 = n7122 | n7683 ;
  assign n15908 = x[82] & n7098 ;
  assign n15909 = n15907 | n15908 ;
  assign n15910 = n7194 | n15909 ;
  assign n28955 = ~n15910 ;
  assign n15911 = x[20] & n28955 ;
  assign n15912 = n28114 & n15910 ;
  assign n15913 = n15911 | n15912 ;
  assign n15914 = n15906 & n15913 ;
  assign n16157 = n15906 | n15913 ;
  assign n28956 = ~n15914 ;
  assign n16459 = n28956 & n16157 ;
  assign n16460 = n16458 & n16459 ;
  assign n16813 = n16458 | n16459 ;
  assign n28957 = ~n16460 ;
  assign n16814 = n28957 & n16813 ;
  assign n8711 = n1239 & n8706 ;
  assign n8661 = x[83] & n8645 ;
  assign n9889 = x[84] & n9278 ;
  assign n16815 = n8661 | n9889 ;
  assign n16816 = x[85] & n8643 ;
  assign n16817 = n16815 | n16816 ;
  assign n16818 = n8711 | n16817 ;
  assign n28958 = ~n16818 ;
  assign n16819 = x[17] & n28958 ;
  assign n16820 = n28039 & n16818 ;
  assign n16821 = n16819 | n16820 ;
  assign n28959 = ~n16821 ;
  assign n16822 = n16814 & n28959 ;
  assign n28960 = ~n16814 ;
  assign n17813 = n28960 & n16821 ;
  assign n17814 = n16822 | n17813 ;
  assign n17815 = n17812 | n17814 ;
  assign n17816 = n17812 & n17814 ;
  assign n28961 = ~n17816 ;
  assign n17844 = n17815 & n28961 ;
  assign n10562 = n1720 & n10542 ;
  assign n10503 = x[86] & n10481 ;
  assign n11915 = x[87] & n11232 ;
  assign n17845 = n10503 | n11915 ;
  assign n17846 = x[88] & n10479 ;
  assign n17847 = n17845 | n17846 ;
  assign n17848 = n10562 | n17847 ;
  assign n28962 = ~n17848 ;
  assign n17849 = x[14] & n28962 ;
  assign n17850 = n27956 & n17848 ;
  assign n17851 = n17849 | n17850 ;
  assign n17852 = n17844 & n17851 ;
  assign n18192 = n17844 | n17851 ;
  assign n28963 = ~n17852 ;
  assign n18708 = n28963 & n18192 ;
  assign n28964 = ~n18191 ;
  assign n18710 = n28964 & n18708 ;
  assign n28965 = ~n18708 ;
  assign n19026 = n18191 & n28965 ;
  assign n19027 = n18710 | n19026 ;
  assign n28966 = ~n19025 ;
  assign n19486 = n28966 & n19027 ;
  assign n28967 = ~n19027 ;
  assign n19487 = n19025 & n28967 ;
  assign n19488 = n19486 | n19487 ;
  assign n28968 = ~n19488 ;
  assign n20060 = n19485 & n28968 ;
  assign n28969 = ~n19485 ;
  assign n20295 = n28969 & n19488 ;
  assign n20296 = n20060 | n20295 ;
  assign n15340 = n2410 & n15308 ;
  assign n15259 = x[92] & n15246 ;
  assign n17298 = x[93] & n16288 ;
  assign n20297 = n15259 | n17298 ;
  assign n20298 = x[94] & n15244 ;
  assign n20299 = n20297 | n20298 ;
  assign n20300 = n15340 | n20299 ;
  assign n28970 = ~n20300 ;
  assign n20301 = x[8] & n28970 ;
  assign n20302 = n27845 & n20300 ;
  assign n20303 = n20301 | n20302 ;
  assign n20304 = n20296 | n20303 ;
  assign n20305 = n20296 & n20303 ;
  assign n28971 = ~n20305 ;
  assign n21241 = n20304 & n28971 ;
  assign n21242 = n21240 & n21241 ;
  assign n21466 = n21240 | n21241 ;
  assign n28972 = ~n21242 ;
  assign n21467 = n28972 & n21466 ;
  assign n21468 = n21465 & n21467 ;
  assign n21952 = n21465 | n21467 ;
  assign n28973 = ~n21468 ;
  assign n21953 = n28973 & n21952 ;
  assign n21954 = n21951 & n21953 ;
  assign n22473 = n21951 | n21953 ;
  assign n28974 = ~n21954 ;
  assign n22474 = n28974 & n22473 ;
  assign n561 = n559 & n560 ;
  assign n562 = n27627 | n561 ;
  assign n25527 = x[99] & x[100] ;
  assign n563 = x[99] | x[100] ;
  assign n28975 = ~n25527 ;
  assign n2463 = n28975 & n563 ;
  assign n2464 = n562 & n2463 ;
  assign n2465 = n562 | n2463 ;
  assign n28976 = ~n2464 ;
  assign n2466 = n28976 & n2465 ;
  assign n19691 = n2466 & n19656 ;
  assign n19754 = x[98] & n19723 ;
  assign n19841 = x[99] & n19829 ;
  assign n22475 = n19754 | n19841 ;
  assign n22476 = x[100] & n19655 ;
  assign n22477 = n22475 | n22476 ;
  assign n22478 = n19691 | n22477 ;
  assign n28977 = ~n22478 ;
  assign n22479 = x[2] & n28977 ;
  assign n22480 = n27790 & n22478 ;
  assign n22481 = n22479 | n22480 ;
  assign n28978 = ~n22481 ;
  assign n22482 = n22474 & n28978 ;
  assign n28979 = ~n22474 ;
  assign n22484 = n28979 & n22481 ;
  assign n22485 = n22482 | n22484 ;
  assign n22995 = n22991 | n22994 ;
  assign n22996 = n22485 & n22995 ;
  assign n27675 = n22485 | n22995 ;
  assign n28980 = ~n22996 ;
  assign n165 = n28980 & n27675 ;
  assign n22483 = n22474 & n22481 ;
  assign n22997 = n22483 | n22996 ;
  assign n21955 = n21468 | n21954 ;
  assign n18449 = n2841 & n18392 ;
  assign n18354 = x[96] & n18329 ;
  assign n18560 = x[97] & n18514 ;
  assign n21446 = n18354 | n18560 ;
  assign n21447 = x[98] & n18327 ;
  assign n21448 = n21446 | n21447 ;
  assign n21449 = n18449 | n21448 ;
  assign n28981 = ~n21449 ;
  assign n21450 = x[5] & n28981 ;
  assign n21451 = n27813 & n21449 ;
  assign n21452 = n21450 | n21451 ;
  assign n15350 = n2152 & n15308 ;
  assign n15271 = x[93] & n15246 ;
  assign n17300 = x[94] & n16288 ;
  assign n20285 = n15271 | n17300 ;
  assign n20286 = x[95] & n15244 ;
  assign n20287 = n20285 | n20286 ;
  assign n20288 = n15350 | n20287 ;
  assign n28982 = ~n20288 ;
  assign n20289 = x[8] & n28982 ;
  assign n20290 = n27845 & n20288 ;
  assign n20291 = n20289 | n20290 ;
  assign n19028 = n19025 & n19027 ;
  assign n19490 = n19485 & n19488 ;
  assign n19491 = n19028 | n19490 ;
  assign n18193 = n18191 & n18192 ;
  assign n18194 = n17852 | n18193 ;
  assign n8763 = n1213 & n8706 ;
  assign n8656 = x[84] & n8645 ;
  assign n9888 = x[85] & n9278 ;
  assign n16800 = n8656 | n9888 ;
  assign n16801 = x[86] & n8643 ;
  assign n16802 = n16800 | n16801 ;
  assign n16803 = n8763 | n16802 ;
  assign n28983 = ~n16803 ;
  assign n16804 = x[17] & n28983 ;
  assign n16805 = n28039 & n16803 ;
  assign n16806 = n16804 | n16805 ;
  assign n5306 = n1270 & n5302 ;
  assign n5268 = x[78] & n5240 ;
  assign n6249 = x[79] & n6179 ;
  assign n14878 = n5268 | n6249 ;
  assign n14879 = x[80] & n5238 ;
  assign n14880 = n14878 | n14879 ;
  assign n14881 = n5306 | n14880 ;
  assign n28984 = ~n14881 ;
  assign n14882 = x[23] & n28984 ;
  assign n14883 = n28221 & n14881 ;
  assign n14884 = n14882 | n14883 ;
  assign n28985 = ~n13364 ;
  assign n13766 = n28985 & n13365 ;
  assign n28986 = ~n13365 ;
  assign n13979 = n13364 & n28986 ;
  assign n13980 = n13766 | n13979 ;
  assign n13989 = n13980 & n13987 ;
  assign n14156 = n13989 | n14155 ;
  assign n1776 = n452 & n1775 ;
  assign n365 = x[75] & n330 ;
  assign n413 = x[76] & n390 ;
  assign n13969 = n365 | n413 ;
  assign n13970 = x[77] & n322 ;
  assign n13971 = n13969 | n13970 ;
  assign n13972 = n1776 | n13971 ;
  assign n28987 = ~n13972 ;
  assign n13973 = x[26] & n28987 ;
  assign n13974 = n28342 & n13972 ;
  assign n13975 = n13973 | n13974 ;
  assign n13367 = n13254 | n13366 ;
  assign n4673 = n2722 & n4632 ;
  assign n4549 = x[72] & n4514 ;
  assign n4616 = x[73] & n4572 ;
  assign n13233 = n4549 | n4616 ;
  assign n13234 = x[74] & n4504 ;
  assign n13235 = n13233 | n13234 ;
  assign n13236 = n4673 | n13235 ;
  assign n28988 = ~n13236 ;
  assign n13237 = x[29] & n28988 ;
  assign n13238 = n28483 & n13236 ;
  assign n13239 = n13237 | n13238 ;
  assign n12381 = n12377 & n12379 ;
  assign n12445 = n12442 & n12444 ;
  assign n12446 = n12381 | n12445 ;
  assign n4792 = n779 & n4790 ;
  assign n714 = x[69] & n663 ;
  assign n769 = x[70] & n720 ;
  assign n12360 = n714 | n769 ;
  assign n12361 = x[71] & n652 ;
  assign n12362 = n12360 | n12361 ;
  assign n12363 = n4792 | n12362 ;
  assign n28989 = ~n12363 ;
  assign n12364 = x[32] & n28989 ;
  assign n12365 = n28658 & n12363 ;
  assign n12366 = n12364 | n12365 ;
  assign n11620 = n11611 & n11618 ;
  assign n11621 = n10992 & n11608 ;
  assign n11622 = n11620 | n11621 ;
  assign n6417 = n4041 & n6408 ;
  assign n3957 = x[66] & n3910 ;
  assign n3980 = x[67] & n3975 ;
  assign n11579 = n3957 | n3980 ;
  assign n11580 = x[68] & n3906 ;
  assign n11581 = n11579 | n11580 ;
  assign n11582 = n6417 | n11581 ;
  assign n11583 = x[35] | n11582 ;
  assign n11584 = x[35] & n11582 ;
  assign n28990 = ~n11584 ;
  assign n11585 = n11583 & n28990 ;
  assign n10993 = x[38] & n28938 ;
  assign n27731 = x[37] & x[38] ;
  assign n3437 = x[37] | x[38] ;
  assign n28991 = ~n27731 ;
  assign n3438 = n28991 & n3437 ;
  assign n3574 = n3436 & n3438 ;
  assign n6446 = n3574 & n6437 ;
  assign n28992 = ~n3438 ;
  assign n3439 = n3436 & n28992 ;
  assign n10994 = x[65] & n3439 ;
  assign n27732 = x[36] & x[37] ;
  assign n3440 = x[36] | x[37] ;
  assign n28993 = ~n27732 ;
  assign n3441 = n28993 & n3440 ;
  assign n28994 = ~n3436 ;
  assign n3508 = n28994 & n3441 ;
  assign n10995 = x[64] & n3508 ;
  assign n10996 = n10994 | n10995 ;
  assign n10997 = n6446 | n10996 ;
  assign n28995 = ~n10997 ;
  assign n10998 = x[38] & n28995 ;
  assign n28996 = ~x[38] ;
  assign n10999 = n28996 & n10997 ;
  assign n11000 = n10998 | n10999 ;
  assign n28997 = ~n11000 ;
  assign n11001 = n10993 & n28997 ;
  assign n28998 = ~n10993 ;
  assign n11586 = n28998 & n11000 ;
  assign n11587 = n11001 | n11586 ;
  assign n11588 = n11585 & n11587 ;
  assign n11623 = n11585 | n11587 ;
  assign n28999 = ~n11588 ;
  assign n11624 = n28999 & n11623 ;
  assign n29000 = ~n11622 ;
  assign n11625 = n29000 & n11624 ;
  assign n29001 = ~n11624 ;
  assign n12367 = n11622 & n29001 ;
  assign n12368 = n11625 | n12367 ;
  assign n12369 = n12366 | n12368 ;
  assign n12370 = n12366 & n12368 ;
  assign n29002 = ~n12370 ;
  assign n12447 = n12369 & n29002 ;
  assign n12448 = n12446 & n12447 ;
  assign n13240 = n12446 | n12447 ;
  assign n29003 = ~n12448 ;
  assign n13241 = n29003 & n13240 ;
  assign n13242 = n13239 & n13241 ;
  assign n13368 = n13239 | n13241 ;
  assign n29004 = ~n13242 ;
  assign n13769 = n29004 & n13368 ;
  assign n29005 = ~n13367 ;
  assign n13771 = n29005 & n13769 ;
  assign n29006 = ~n13769 ;
  assign n13976 = n13367 & n29006 ;
  assign n13977 = n13771 | n13976 ;
  assign n13978 = n13975 & n13977 ;
  assign n14157 = n13975 | n13977 ;
  assign n29007 = ~n13978 ;
  assign n14158 = n29007 & n14157 ;
  assign n14159 = n14156 & n14158 ;
  assign n14885 = n14156 | n14158 ;
  assign n29008 = ~n14159 ;
  assign n14886 = n29008 & n14885 ;
  assign n29009 = ~n14884 ;
  assign n14888 = n29009 & n14886 ;
  assign n29010 = ~n14886 ;
  assign n14889 = n14884 & n29010 ;
  assign n14890 = n14888 | n14889 ;
  assign n13988 = n13980 | n13987 ;
  assign n29011 = ~n13989 ;
  assign n14702 = n13988 & n29011 ;
  assign n29012 = ~n14153 ;
  assign n14703 = n29012 & n14702 ;
  assign n29013 = ~n14702 ;
  assign n14898 = n14153 & n29013 ;
  assign n14899 = n14703 | n14898 ;
  assign n14900 = n14897 & n14899 ;
  assign n15091 = n14910 & n15089 ;
  assign n15092 = n14911 | n15091 ;
  assign n15094 = n14897 & n15093 ;
  assign n15096 = n14897 | n15093 ;
  assign n29014 = ~n15094 ;
  assign n15097 = n29014 & n15096 ;
  assign n15098 = n15092 & n15097 ;
  assign n15099 = n14900 | n15098 ;
  assign n15100 = n14890 | n15099 ;
  assign n15101 = n14890 & n15099 ;
  assign n29015 = ~n15101 ;
  assign n15891 = n15100 & n29015 ;
  assign n7172 = n1057 & n7162 ;
  assign n7136 = x[81] & n7100 ;
  assign n7712 = x[82] & n7647 ;
  assign n15892 = n7136 | n7712 ;
  assign n15893 = x[83] & n7098 ;
  assign n15894 = n15892 | n15893 ;
  assign n15895 = n7172 | n15894 ;
  assign n29016 = ~n15895 ;
  assign n15896 = x[20] & n29016 ;
  assign n15897 = n28114 & n15895 ;
  assign n15898 = n15896 | n15897 ;
  assign n29017 = ~n15898 ;
  assign n15899 = n15891 & n29017 ;
  assign n29018 = ~n15891 ;
  assign n16416 = n29018 & n15898 ;
  assign n16417 = n15899 | n16416 ;
  assign n16461 = n15914 | n16460 ;
  assign n16463 = n16417 | n16461 ;
  assign n16464 = n16417 & n16461 ;
  assign n29019 = ~n16464 ;
  assign n16809 = n16463 & n29019 ;
  assign n29020 = ~n16806 ;
  assign n16810 = n29020 & n16809 ;
  assign n29021 = ~n16809 ;
  assign n16811 = n16806 & n29021 ;
  assign n16812 = n16810 | n16811 ;
  assign n16823 = n16814 & n16821 ;
  assign n17114 = n16814 | n16821 ;
  assign n29022 = ~n16823 ;
  assign n17115 = n29022 & n17114 ;
  assign n17116 = n17113 & n17115 ;
  assign n17117 = n16823 | n17116 ;
  assign n17118 = n16812 | n17117 ;
  assign n17119 = n16812 & n17117 ;
  assign n29023 = ~n17119 ;
  assign n17835 = n17118 & n29023 ;
  assign n10563 = n1453 & n10542 ;
  assign n10504 = x[87] & n10481 ;
  assign n11906 = x[88] & n11232 ;
  assign n17836 = n10504 | n11906 ;
  assign n17837 = x[89] & n10479 ;
  assign n17838 = n17836 | n17837 ;
  assign n17839 = n10563 | n17838 ;
  assign n29024 = ~n17839 ;
  assign n17840 = x[14] & n29024 ;
  assign n17841 = n27956 & n17839 ;
  assign n17842 = n17840 | n17841 ;
  assign n17843 = n17835 & n17842 ;
  assign n14887 = n14884 & n14886 ;
  assign n15736 = n14884 | n14886 ;
  assign n29025 = ~n14887 ;
  assign n15737 = n29025 & n15736 ;
  assign n29026 = ~n15099 ;
  assign n15738 = n29026 & n15737 ;
  assign n29027 = ~n15737 ;
  assign n15901 = n15099 & n29027 ;
  assign n15902 = n15738 | n15901 ;
  assign n15903 = n15898 | n15902 ;
  assign n15904 = n15898 & n15902 ;
  assign n29028 = ~n15904 ;
  assign n15905 = n15903 & n29028 ;
  assign n29029 = ~n16461 ;
  assign n16462 = n15905 & n29029 ;
  assign n29030 = ~n15905 ;
  assign n16798 = n29030 & n16461 ;
  assign n16799 = n16462 | n16798 ;
  assign n16807 = n16799 | n16806 ;
  assign n16808 = n16799 & n16806 ;
  assign n29031 = ~n16808 ;
  assign n17753 = n16807 & n29031 ;
  assign n29032 = ~n17117 ;
  assign n17754 = n29032 & n17753 ;
  assign n29033 = ~n17753 ;
  assign n18702 = n17117 & n29033 ;
  assign n18703 = n17754 | n18702 ;
  assign n18712 = n17842 | n18703 ;
  assign n29034 = ~n17843 ;
  assign n19006 = n29034 & n18712 ;
  assign n29035 = ~n19006 ;
  assign n19007 = n18194 & n29035 ;
  assign n18704 = n17842 & n18703 ;
  assign n18705 = n17856 | n17863 ;
  assign n18706 = n18187 & n18705 ;
  assign n18707 = n17865 | n18706 ;
  assign n18709 = n18707 & n18708 ;
  assign n18711 = n17852 | n18709 ;
  assign n18713 = n18711 & n18712 ;
  assign n18714 = n18704 | n18713 ;
  assign n29036 = ~n18714 ;
  assign n19008 = n18712 & n29036 ;
  assign n19009 = n19007 | n19008 ;
  assign n12717 = n1841 & n12695 ;
  assign n12652 = x[90] & n12633 ;
  assign n14367 = x[91] & n13533 ;
  assign n19010 = n12652 | n14367 ;
  assign n19011 = x[92] & n12631 ;
  assign n19012 = n19010 | n19011 ;
  assign n19013 = n12717 | n19012 ;
  assign n29037 = ~n19013 ;
  assign n19014 = x[11] & n29037 ;
  assign n19015 = n27892 & n19013 ;
  assign n19016 = n19014 | n19015 ;
  assign n29038 = ~n19016 ;
  assign n19017 = n19009 & n29038 ;
  assign n29039 = ~n19009 ;
  assign n19492 = n29039 & n19016 ;
  assign n19493 = n19017 | n19492 ;
  assign n19494 = n19491 & n19493 ;
  assign n20292 = n19491 | n19493 ;
  assign n29040 = ~n19494 ;
  assign n20293 = n29040 & n20292 ;
  assign n20294 = n20291 & n20293 ;
  assign n20835 = n20291 | n20293 ;
  assign n29041 = ~n20294 ;
  assign n20836 = n29041 & n20835 ;
  assign n19489 = n19485 | n19488 ;
  assign n29042 = ~n19490 ;
  assign n20831 = n19489 & n29042 ;
  assign n21122 = n20303 & n20831 ;
  assign n21243 = n21122 | n21242 ;
  assign n29043 = ~n21243 ;
  assign n21244 = n20836 & n29043 ;
  assign n29044 = ~n20836 ;
  assign n21453 = n29044 & n21243 ;
  assign n21454 = n21244 | n21453 ;
  assign n21455 = n21452 & n21454 ;
  assign n22103 = n21452 | n21454 ;
  assign n29045 = ~n21455 ;
  assign n22104 = n29045 & n22103 ;
  assign n29046 = ~n21955 ;
  assign n22105 = n29046 & n22104 ;
  assign n29047 = ~n22104 ;
  assign n22462 = n21955 & n29047 ;
  assign n22463 = n22105 | n22462 ;
  assign n564 = n562 & n563 ;
  assign n565 = n25527 | n564 ;
  assign n27625 = x[100] & x[101] ;
  assign n566 = x[100] | x[101] ;
  assign n29048 = ~n27625 ;
  assign n2974 = n29048 & n566 ;
  assign n29049 = ~n565 ;
  assign n2975 = n29049 & n2974 ;
  assign n29050 = ~n2974 ;
  assign n2976 = n565 & n29050 ;
  assign n2977 = n2975 | n2976 ;
  assign n19717 = n2977 & n19656 ;
  assign n19783 = x[99] & n19723 ;
  assign n19888 = x[100] & n19829 ;
  assign n22464 = n19783 | n19888 ;
  assign n22465 = x[101] & n19655 ;
  assign n22466 = n22464 | n22465 ;
  assign n22467 = n19717 | n22466 ;
  assign n29051 = ~n22467 ;
  assign n22468 = x[2] & n29051 ;
  assign n22469 = n27790 & n22467 ;
  assign n22470 = n22468 | n22469 ;
  assign n22471 = n22463 | n22470 ;
  assign n22472 = n22463 & n22470 ;
  assign n29052 = ~n22472 ;
  assign n22998 = n22471 & n29052 ;
  assign n22999 = n22997 | n22998 ;
  assign n23000 = n22997 & n22998 ;
  assign n29053 = ~n23000 ;
  assign n166 = n22999 & n29053 ;
  assign n567 = n565 & n566 ;
  assign n568 = n27625 | n567 ;
  assign n25376 = x[101] & x[102] ;
  assign n569 = x[101] | x[102] ;
  assign n29054 = ~n25376 ;
  assign n2864 = n29054 & n569 ;
  assign n2865 = n568 & n2864 ;
  assign n2866 = n568 | n2864 ;
  assign n29055 = ~n2865 ;
  assign n2867 = n29055 & n2866 ;
  assign n19713 = n2867 & n19656 ;
  assign n19763 = x[100] & n19723 ;
  assign n19887 = x[101] & n19829 ;
  assign n22450 = n19763 | n19887 ;
  assign n22451 = x[102] & n19655 ;
  assign n22452 = n22450 | n22451 ;
  assign n22453 = n19713 | n22452 ;
  assign n22454 = x[2] | n22453 ;
  assign n22455 = x[2] & n22453 ;
  assign n29056 = ~n22455 ;
  assign n22456 = n22454 & n29056 ;
  assign n29057 = ~n21452 ;
  assign n21456 = n29057 & n21454 ;
  assign n29058 = ~n21454 ;
  assign n21457 = n21452 & n29058 ;
  assign n21458 = n21456 | n21457 ;
  assign n21956 = n21458 & n21955 ;
  assign n21957 = n21455 | n21956 ;
  assign n18427 = n2313 & n18392 ;
  assign n18352 = x[97] & n18329 ;
  assign n18568 = x[98] & n18514 ;
  assign n21436 = n18352 | n18568 ;
  assign n21437 = x[99] & n18327 ;
  assign n21438 = n21436 | n21437 ;
  assign n21439 = n18427 | n21438 ;
  assign n29059 = ~n21439 ;
  assign n21440 = x[5] & n29059 ;
  assign n21441 = n27813 & n21439 ;
  assign n21442 = n21440 | n21441 ;
  assign n20828 = n20422 | n20827 ;
  assign n20829 = n20318 & n20828 ;
  assign n20830 = n20315 | n20829 ;
  assign n20832 = n20303 | n20831 ;
  assign n20833 = n20830 & n20832 ;
  assign n20834 = n20305 | n20833 ;
  assign n20837 = n20834 & n20836 ;
  assign n20838 = n20294 | n20837 ;
  assign n15359 = n2000 & n15308 ;
  assign n15260 = x[94] & n15246 ;
  assign n17279 = x[95] & n16288 ;
  assign n20275 = n15260 | n17279 ;
  assign n20276 = x[96] & n15244 ;
  assign n20277 = n20275 | n20276 ;
  assign n20278 = n15359 | n20277 ;
  assign n29060 = ~n20278 ;
  assign n20279 = x[8] & n29060 ;
  assign n20280 = n27845 & n20278 ;
  assign n20281 = n20279 | n20280 ;
  assign n19018 = n19009 & n19016 ;
  assign n19495 = n19018 | n19494 ;
  assign n12719 = n1685 & n12695 ;
  assign n12653 = x[91] & n12633 ;
  assign n14386 = x[92] & n13533 ;
  assign n18996 = n12653 | n14386 ;
  assign n18997 = x[93] & n12631 ;
  assign n18998 = n18996 | n18997 ;
  assign n18999 = n12719 | n18998 ;
  assign n29061 = ~n18999 ;
  assign n19000 = x[11] & n29061 ;
  assign n19001 = n27892 & n18999 ;
  assign n19002 = n19000 | n19001 ;
  assign n18195 = n17835 | n17842 ;
  assign n18196 = n18194 & n18195 ;
  assign n18197 = n17843 | n18196 ;
  assign n17120 = n16808 | n17119 ;
  assign n7173 = n1293 & n7162 ;
  assign n7127 = x[82] & n7100 ;
  assign n7685 = x[83] & n7647 ;
  assign n15878 = n7127 | n7685 ;
  assign n15879 = x[84] & n7098 ;
  assign n15880 = n15878 | n15879 ;
  assign n15881 = n7173 | n15880 ;
  assign n29062 = ~n15881 ;
  assign n15882 = x[20] & n29062 ;
  assign n15883 = n28114 & n15881 ;
  assign n15884 = n15882 | n15883 ;
  assign n5308 = n1029 & n5302 ;
  assign n5272 = x[79] & n5240 ;
  assign n6229 = x[80] & n6179 ;
  assign n14865 = n5272 | n6229 ;
  assign n14866 = x[81] & n5238 ;
  assign n14867 = n14865 | n14866 ;
  assign n14868 = n5308 | n14867 ;
  assign n29063 = ~n14868 ;
  assign n14869 = x[23] & n29063 ;
  assign n14870 = n28221 & n14868 ;
  assign n14871 = n14869 | n14870 ;
  assign n14160 = n13978 | n14159 ;
  assign n4634 = n3289 & n4632 ;
  assign n4521 = x[73] & n4514 ;
  assign n4621 = x[74] & n4572 ;
  assign n13222 = n4521 | n4621 ;
  assign n13223 = x[75] & n4504 ;
  assign n13224 = n13222 | n13223 ;
  assign n13225 = n4634 | n13224 ;
  assign n29064 = ~n13225 ;
  assign n13226 = x[29] & n29064 ;
  assign n13227 = n28483 & n13225 ;
  assign n13228 = n13226 | n13227 ;
  assign n12449 = n12370 | n12448 ;
  assign n11626 = n11622 & n11624 ;
  assign n11627 = n11588 | n11626 ;
  assign n11002 = n10993 & n11000 ;
  assign n6470 = n3574 & n6466 ;
  assign n3442 = n28994 & n3438 ;
  assign n29065 = ~n3441 ;
  assign n3443 = n29065 & n3442 ;
  assign n3477 = x[64] & n3443 ;
  assign n3555 = x[65] & n3508 ;
  assign n11003 = n3477 | n3555 ;
  assign n11004 = x[66] & n3439 ;
  assign n11005 = n11003 | n11004 ;
  assign n11006 = n6470 | n11005 ;
  assign n29066 = ~n11006 ;
  assign n11007 = x[38] & n29066 ;
  assign n11008 = n28996 & n11006 ;
  assign n11009 = n11007 | n11008 ;
  assign n29067 = ~n11009 ;
  assign n11010 = n11002 & n29067 ;
  assign n29068 = ~n11002 ;
  assign n11568 = n29068 & n11009 ;
  assign n11569 = n11010 | n11568 ;
  assign n6380 = n4041 & n6379 ;
  assign n3916 = x[67] & n3910 ;
  assign n3981 = x[68] & n3975 ;
  assign n11570 = n3916 | n3981 ;
  assign n11571 = x[69] & n3906 ;
  assign n11572 = n11570 | n11571 ;
  assign n11573 = n6380 | n11572 ;
  assign n29069 = ~n11573 ;
  assign n11574 = x[35] & n29069 ;
  assign n11575 = n28822 & n11573 ;
  assign n11576 = n11574 | n11575 ;
  assign n29070 = ~n11576 ;
  assign n11577 = n11569 & n29070 ;
  assign n29071 = ~n11569 ;
  assign n11628 = n29071 & n11576 ;
  assign n11629 = n11577 | n11628 ;
  assign n11630 = n11627 & n11629 ;
  assign n12349 = n11627 | n11629 ;
  assign n29072 = ~n11630 ;
  assign n12350 = n29072 & n12349 ;
  assign n3702 = n779 & n3701 ;
  assign n706 = x[70] & n663 ;
  assign n757 = x[71] & n720 ;
  assign n12351 = n706 | n757 ;
  assign n12352 = x[72] & n652 ;
  assign n12353 = n12351 | n12352 ;
  assign n12354 = n3702 | n12353 ;
  assign n29073 = ~n12354 ;
  assign n12355 = x[32] & n29073 ;
  assign n12356 = n28658 & n12354 ;
  assign n12357 = n12355 | n12356 ;
  assign n12358 = n12350 | n12357 ;
  assign n12359 = n12350 & n12357 ;
  assign n29074 = ~n12359 ;
  assign n12450 = n12358 & n29074 ;
  assign n29075 = ~n12449 ;
  assign n12451 = n29075 & n12450 ;
  assign n29076 = ~n12450 ;
  assign n13229 = n12449 & n29076 ;
  assign n13230 = n12451 | n13229 ;
  assign n29077 = ~n13228 ;
  assign n13231 = n29077 & n13230 ;
  assign n29078 = ~n13230 ;
  assign n13371 = n13228 & n29078 ;
  assign n13372 = n13231 | n13371 ;
  assign n13767 = n13253 & n13364 ;
  assign n13768 = n13254 | n13767 ;
  assign n13770 = n13768 & n13769 ;
  assign n13772 = n13242 | n13770 ;
  assign n13773 = n13372 | n13772 ;
  assign n13774 = n13372 & n13772 ;
  assign n29079 = ~n13774 ;
  assign n13959 = n13773 & n29079 ;
  assign n2087 = n452 & n2084 ;
  assign n355 = x[76] & n330 ;
  assign n442 = x[77] & n390 ;
  assign n13960 = n355 | n442 ;
  assign n13961 = x[78] & n322 ;
  assign n13962 = n13960 | n13961 ;
  assign n13963 = n2087 | n13962 ;
  assign n29080 = ~n13963 ;
  assign n13964 = x[26] & n29080 ;
  assign n13965 = n28342 & n13963 ;
  assign n13966 = n13964 | n13965 ;
  assign n13967 = n13959 | n13966 ;
  assign n13968 = n13959 & n13966 ;
  assign n29081 = ~n13968 ;
  assign n14721 = n13967 & n29081 ;
  assign n29082 = ~n14160 ;
  assign n14723 = n29082 & n14721 ;
  assign n29083 = ~n14721 ;
  assign n14872 = n14160 & n29083 ;
  assign n14873 = n14723 | n14872 ;
  assign n29084 = ~n14871 ;
  assign n14875 = n29084 & n14873 ;
  assign n29085 = ~n14873 ;
  assign n15734 = n14871 & n29085 ;
  assign n15735 = n14875 | n15734 ;
  assign n15777 = n14900 | n15776 ;
  assign n15778 = n15737 & n15777 ;
  assign n15779 = n14887 | n15778 ;
  assign n15781 = n15735 | n15779 ;
  assign n15782 = n15735 & n15779 ;
  assign n29086 = ~n15782 ;
  assign n15887 = n15781 & n29086 ;
  assign n29087 = ~n15884 ;
  assign n15888 = n29087 & n15887 ;
  assign n29088 = ~n15887 ;
  assign n15889 = n15884 & n29088 ;
  assign n15890 = n15888 | n15889 ;
  assign n15900 = n15891 & n15898 ;
  assign n16154 = n15938 | n16153 ;
  assign n16155 = n15927 & n16154 ;
  assign n16156 = n15924 | n16155 ;
  assign n16158 = n16156 & n16157 ;
  assign n16159 = n15914 | n16158 ;
  assign n16160 = n15905 & n16159 ;
  assign n16161 = n15900 | n16160 ;
  assign n16162 = n15890 | n16161 ;
  assign n16163 = n15890 & n16161 ;
  assign n29089 = ~n16163 ;
  assign n16789 = n16162 & n29089 ;
  assign n8720 = n1522 & n8706 ;
  assign n8658 = x[85] & n8645 ;
  assign n9887 = x[86] & n9278 ;
  assign n16790 = n8658 | n9887 ;
  assign n16791 = x[87] & n8643 ;
  assign n16792 = n16790 | n16791 ;
  assign n16793 = n8720 | n16792 ;
  assign n29090 = ~n16793 ;
  assign n16794 = x[17] & n29090 ;
  assign n16795 = n28039 & n16793 ;
  assign n16796 = n16794 | n16795 ;
  assign n16797 = n16789 & n16796 ;
  assign n14874 = n14871 & n14873 ;
  assign n14876 = n14871 | n14873 ;
  assign n29091 = ~n14874 ;
  assign n14877 = n29091 & n14876 ;
  assign n29092 = ~n15779 ;
  assign n15780 = n14877 & n29092 ;
  assign n29093 = ~n14877 ;
  assign n15876 = n29093 & n15779 ;
  assign n15877 = n15780 | n15876 ;
  assign n15885 = n15877 | n15884 ;
  assign n15886 = n15877 & n15884 ;
  assign n29094 = ~n15886 ;
  assign n16414 = n15885 & n29094 ;
  assign n29095 = ~n16161 ;
  assign n16415 = n29095 & n16414 ;
  assign n29096 = ~n16414 ;
  assign n17748 = n16161 & n29096 ;
  assign n17749 = n16415 | n17748 ;
  assign n17750 = n16796 | n17749 ;
  assign n29097 = ~n16797 ;
  assign n17822 = n29097 & n17750 ;
  assign n29098 = ~n17822 ;
  assign n17823 = n17120 & n29098 ;
  assign n17751 = n16796 & n17749 ;
  assign n17752 = n16806 & n16809 ;
  assign n17817 = n16823 | n17816 ;
  assign n17818 = n17753 & n17817 ;
  assign n17819 = n17752 | n17818 ;
  assign n17820 = n17750 & n17819 ;
  assign n17821 = n17751 | n17820 ;
  assign n29099 = ~n17821 ;
  assign n17824 = n17750 & n29099 ;
  assign n17825 = n17823 | n17824 ;
  assign n10578 = n1482 & n10542 ;
  assign n10526 = x[88] & n10481 ;
  assign n11913 = x[89] & n11232 ;
  assign n17826 = n10526 | n11913 ;
  assign n17827 = x[90] & n10479 ;
  assign n17828 = n17826 | n17827 ;
  assign n17829 = n10578 | n17828 ;
  assign n29100 = ~n17829 ;
  assign n17830 = x[14] & n29100 ;
  assign n17831 = n27956 & n17829 ;
  assign n17832 = n17830 | n17831 ;
  assign n29101 = ~n17832 ;
  assign n17833 = n17825 & n29101 ;
  assign n29102 = ~n17825 ;
  assign n18715 = n29102 & n17832 ;
  assign n18716 = n17833 | n18715 ;
  assign n29103 = ~n18197 ;
  assign n18718 = n29103 & n18716 ;
  assign n29104 = ~n18716 ;
  assign n19003 = n18197 & n29104 ;
  assign n19004 = n18718 | n19003 ;
  assign n19005 = n19002 & n19004 ;
  assign n19496 = n19002 | n19004 ;
  assign n29105 = ~n19005 ;
  assign n20068 = n29105 & n19496 ;
  assign n29106 = ~n19495 ;
  assign n20070 = n29106 & n20068 ;
  assign n29107 = ~n20068 ;
  assign n20282 = n19495 & n29107 ;
  assign n20283 = n20070 | n20282 ;
  assign n20284 = n20281 & n20283 ;
  assign n20839 = n20281 | n20283 ;
  assign n29108 = ~n20284 ;
  assign n21247 = n29108 & n20839 ;
  assign n29109 = ~n20838 ;
  assign n21249 = n29109 & n21247 ;
  assign n29110 = ~n21247 ;
  assign n21443 = n20838 & n29110 ;
  assign n21444 = n21249 | n21443 ;
  assign n21445 = n21442 & n21444 ;
  assign n21958 = n21442 | n21444 ;
  assign n29111 = ~n21445 ;
  assign n21959 = n29111 & n21958 ;
  assign n21960 = n21957 & n21959 ;
  assign n22457 = n21957 | n21959 ;
  assign n29112 = ~n21960 ;
  assign n22458 = n29112 & n22457 ;
  assign n22459 = n22456 & n22458 ;
  assign n22460 = n22456 | n22458 ;
  assign n29113 = ~n22459 ;
  assign n22461 = n29113 & n22460 ;
  assign n23001 = n22472 | n23000 ;
  assign n23002 = n22461 & n23001 ;
  assign n27678 = n22461 | n23001 ;
  assign n29114 = ~n23002 ;
  assign n167 = n29114 & n27678 ;
  assign n570 = n568 & n569 ;
  assign n571 = n25376 | n570 ;
  assign n27624 = x[102] & x[103] ;
  assign n572 = x[102] | x[103] ;
  assign n29115 = ~n27624 ;
  assign n2623 = n29115 & n572 ;
  assign n29116 = ~n571 ;
  assign n2624 = n29116 & n2623 ;
  assign n29117 = ~n2623 ;
  assign n2625 = n571 & n29117 ;
  assign n2626 = n2624 | n2625 ;
  assign n19700 = n2626 & n19656 ;
  assign n19764 = x[101] & n19723 ;
  assign n19885 = x[102] & n19829 ;
  assign n22437 = n19764 | n19885 ;
  assign n22438 = x[103] & n19655 ;
  assign n22439 = n22437 | n22438 ;
  assign n22440 = n19700 | n22439 ;
  assign n29118 = ~n22440 ;
  assign n22441 = x[2] & n29118 ;
  assign n22442 = n27790 & n22440 ;
  assign n22443 = n22441 | n22442 ;
  assign n21961 = n21445 | n21960 ;
  assign n21245 = n20835 & n21243 ;
  assign n21246 = n20294 | n21245 ;
  assign n21248 = n21246 & n21247 ;
  assign n21250 = n20284 | n21248 ;
  assign n15360 = n2438 & n15308 ;
  assign n15261 = x[95] & n15246 ;
  assign n17327 = x[96] & n16288 ;
  assign n20265 = n15261 | n17327 ;
  assign n20266 = x[97] & n15244 ;
  assign n20267 = n20265 | n20266 ;
  assign n20268 = n15360 | n20267 ;
  assign n29119 = ~n20268 ;
  assign n20269 = x[8] & n29119 ;
  assign n20270 = n27845 & n20268 ;
  assign n20271 = n20269 | n20270 ;
  assign n17834 = n17825 & n17832 ;
  assign n18717 = n18714 & n18716 ;
  assign n18719 = n17834 | n18717 ;
  assign n10600 = n2046 & n10542 ;
  assign n10506 = x[89] & n10481 ;
  assign n11912 = x[90] & n11232 ;
  assign n17738 = n10506 | n11912 ;
  assign n17739 = x[91] & n10479 ;
  assign n17740 = n17738 | n17739 ;
  assign n17741 = n10600 | n17740 ;
  assign n29120 = ~n17741 ;
  assign n17742 = x[14] & n29120 ;
  assign n17743 = n27956 & n17741 ;
  assign n17744 = n17742 | n17743 ;
  assign n17121 = n16789 | n16796 ;
  assign n17122 = n17120 & n17121 ;
  assign n17123 = n16797 | n17122 ;
  assign n15783 = n14874 | n15782 ;
  assign n14701 = n13987 & n13991 ;
  assign n14706 = n14138 & n14704 ;
  assign n14707 = n14041 | n14706 ;
  assign n14708 = n14028 & n14707 ;
  assign n14709 = n14029 | n14708 ;
  assign n14710 = n14017 & n14709 ;
  assign n14711 = n14015 | n14710 ;
  assign n14715 = n14711 & n14713 ;
  assign n14716 = n14004 | n14715 ;
  assign n14717 = n14702 & n14716 ;
  assign n14718 = n14701 | n14717 ;
  assign n14719 = n14157 & n14718 ;
  assign n14720 = n13978 | n14719 ;
  assign n14722 = n14720 & n14721 ;
  assign n14724 = n13968 | n14722 ;
  assign n1742 = n452 & n1741 ;
  assign n345 = x[77] & n330 ;
  assign n399 = x[78] & n390 ;
  assign n13949 = n345 | n399 ;
  assign n13950 = x[79] & n322 ;
  assign n13951 = n13949 | n13950 ;
  assign n13952 = n1742 | n13951 ;
  assign n29121 = ~n13952 ;
  assign n13953 = x[26] & n29121 ;
  assign n13954 = n28342 & n13952 ;
  assign n13955 = n13953 | n13954 ;
  assign n5983 = n4041 & n5976 ;
  assign n3917 = x[68] & n3910 ;
  assign n3983 = x[69] & n3975 ;
  assign n11556 = n3917 | n3983 ;
  assign n11557 = x[70] & n3906 ;
  assign n11558 = n11556 | n11557 ;
  assign n11559 = n5983 | n11558 ;
  assign n29122 = ~n11559 ;
  assign n11560 = x[35] & n29122 ;
  assign n11561 = n28822 & n11559 ;
  assign n11562 = n11560 | n11561 ;
  assign n27722 = x[38] & x[39] ;
  assign n3023 = x[38] | x[39] ;
  assign n29123 = ~n27722 ;
  assign n3024 = n29123 & n3023 ;
  assign n10239 = x[64] & n3024 ;
  assign n11011 = n11002 & n11009 ;
  assign n11012 = n10239 & n11011 ;
  assign n11013 = n10239 | n11011 ;
  assign n29124 = ~n11012 ;
  assign n11014 = n29124 & n11013 ;
  assign n6500 = n3574 & n6494 ;
  assign n3450 = x[65] & n3443 ;
  assign n3534 = x[66] & n3508 ;
  assign n11015 = n3450 | n3534 ;
  assign n11016 = x[67] & n3439 ;
  assign n11017 = n11015 | n11016 ;
  assign n11018 = n6500 | n11017 ;
  assign n29125 = ~n11018 ;
  assign n11019 = x[38] & n29125 ;
  assign n11020 = n28996 & n11018 ;
  assign n11021 = n11019 | n11020 ;
  assign n29126 = ~n11021 ;
  assign n11022 = n11014 & n29126 ;
  assign n29127 = ~n11014 ;
  assign n11563 = n29127 & n11021 ;
  assign n11564 = n11022 | n11563 ;
  assign n11565 = n11562 & n11564 ;
  assign n11566 = n11562 | n11564 ;
  assign n29128 = ~n11565 ;
  assign n11567 = n29128 & n11566 ;
  assign n11578 = n11569 & n11576 ;
  assign n11631 = n11578 | n11630 ;
  assign n29129 = ~n11631 ;
  assign n11632 = n11567 & n29129 ;
  assign n29130 = ~n11567 ;
  assign n12336 = n29130 & n11631 ;
  assign n12337 = n11632 | n12336 ;
  assign n3734 = n779 & n3733 ;
  assign n691 = x[71] & n663 ;
  assign n735 = x[72] & n720 ;
  assign n12338 = n691 | n735 ;
  assign n12339 = x[73] & n652 ;
  assign n12340 = n12338 | n12339 ;
  assign n12341 = n3734 | n12340 ;
  assign n29131 = ~n12341 ;
  assign n12342 = x[32] & n29131 ;
  assign n12343 = n28658 & n12341 ;
  assign n12344 = n12342 | n12343 ;
  assign n29132 = ~n12344 ;
  assign n12345 = n12337 & n29132 ;
  assign n29133 = ~n12337 ;
  assign n12347 = n29133 & n12344 ;
  assign n12348 = n12345 | n12347 ;
  assign n12452 = n12449 & n12450 ;
  assign n12453 = n12359 | n12452 ;
  assign n12454 = n12348 | n12453 ;
  assign n12455 = n12348 & n12453 ;
  assign n29134 = ~n12455 ;
  assign n13210 = n12454 & n29134 ;
  assign n4650 = n2750 & n4632 ;
  assign n4563 = x[74] & n4514 ;
  assign n4600 = x[75] & n4572 ;
  assign n13211 = n4563 | n4600 ;
  assign n13212 = x[76] & n4504 ;
  assign n13213 = n13211 | n13212 ;
  assign n13214 = n4650 | n13213 ;
  assign n29135 = ~n13214 ;
  assign n13215 = x[29] & n29135 ;
  assign n13216 = n28483 & n13214 ;
  assign n13217 = n13215 | n13216 ;
  assign n29136 = ~n13217 ;
  assign n13218 = n13210 & n29136 ;
  assign n29137 = ~n13210 ;
  assign n13220 = n29137 & n13217 ;
  assign n13221 = n13218 | n13220 ;
  assign n13232 = n13228 & n13230 ;
  assign n13369 = n13367 & n13368 ;
  assign n13370 = n13242 | n13369 ;
  assign n13373 = n13370 & n13372 ;
  assign n13374 = n13232 | n13373 ;
  assign n13376 = n13221 | n13374 ;
  assign n13377 = n13221 & n13374 ;
  assign n29138 = ~n13377 ;
  assign n14163 = n13376 & n29138 ;
  assign n29139 = ~n13955 ;
  assign n14165 = n29139 & n14163 ;
  assign n29140 = ~n14163 ;
  assign n14725 = n13955 & n29140 ;
  assign n14726 = n14165 | n14725 ;
  assign n14727 = n14724 | n14726 ;
  assign n14728 = n14724 & n14726 ;
  assign n29141 = ~n14728 ;
  assign n14855 = n14727 & n29141 ;
  assign n5325 = n1003 & n5302 ;
  assign n5250 = x[80] & n5240 ;
  assign n6231 = x[81] & n6179 ;
  assign n14856 = n5250 | n6231 ;
  assign n14857 = x[82] & n5238 ;
  assign n14858 = n14856 | n14857 ;
  assign n14859 = n5325 | n14858 ;
  assign n29142 = ~n14859 ;
  assign n14860 = x[23] & n29142 ;
  assign n14861 = n28221 & n14859 ;
  assign n14862 = n14860 | n14861 ;
  assign n14863 = n14855 | n14862 ;
  assign n14864 = n14855 & n14862 ;
  assign n29143 = ~n14864 ;
  assign n15784 = n14863 & n29143 ;
  assign n15785 = n15783 & n15784 ;
  assign n15863 = n15783 | n15784 ;
  assign n29144 = ~n15785 ;
  assign n15864 = n29144 & n15863 ;
  assign n7186 = n1239 & n7162 ;
  assign n7131 = x[83] & n7100 ;
  assign n7702 = x[84] & n7647 ;
  assign n15865 = n7131 | n7702 ;
  assign n15866 = x[85] & n7098 ;
  assign n15867 = n15865 | n15866 ;
  assign n15868 = n7186 | n15867 ;
  assign n29145 = ~n15868 ;
  assign n15869 = x[20] & n29145 ;
  assign n15870 = n28114 & n15868 ;
  assign n15871 = n15869 | n15870 ;
  assign n15873 = n15864 & n15871 ;
  assign n15874 = n15864 | n15871 ;
  assign n29146 = ~n15873 ;
  assign n15875 = n29146 & n15874 ;
  assign n16413 = n15884 & n15887 ;
  assign n16465 = n15904 | n16464 ;
  assign n16466 = n16414 & n16465 ;
  assign n16467 = n16413 | n16466 ;
  assign n29147 = ~n16467 ;
  assign n16468 = n15875 & n29147 ;
  assign n29148 = ~n15875 ;
  assign n16778 = n29148 & n16467 ;
  assign n16779 = n16468 | n16778 ;
  assign n8739 = n1720 & n8706 ;
  assign n8659 = x[86] & n8645 ;
  assign n9845 = x[87] & n9278 ;
  assign n16780 = n8659 | n9845 ;
  assign n16781 = x[88] & n8643 ;
  assign n16782 = n16780 | n16781 ;
  assign n16783 = n8739 | n16782 ;
  assign n29149 = ~n16783 ;
  assign n16784 = x[17] & n29149 ;
  assign n16785 = n28039 & n16783 ;
  assign n16786 = n16784 | n16785 ;
  assign n16787 = n16779 | n16786 ;
  assign n16788 = n16779 & n16786 ;
  assign n29150 = ~n16788 ;
  assign n17124 = n16787 & n29150 ;
  assign n29151 = ~n17123 ;
  assign n17125 = n29151 & n17124 ;
  assign n29152 = ~n17124 ;
  assign n17745 = n17123 & n29152 ;
  assign n17746 = n17125 | n17745 ;
  assign n29153 = ~n17744 ;
  assign n18201 = n29153 & n17746 ;
  assign n29154 = ~n17746 ;
  assign n18720 = n17744 & n29154 ;
  assign n18721 = n18201 | n18720 ;
  assign n18722 = n18719 | n18721 ;
  assign n18723 = n18719 & n18721 ;
  assign n29155 = ~n18723 ;
  assign n18987 = n18722 & n29155 ;
  assign n12736 = n2410 & n12695 ;
  assign n12656 = x[92] & n12633 ;
  assign n14351 = x[93] & n13533 ;
  assign n18988 = n12656 | n14351 ;
  assign n18989 = x[94] & n12631 ;
  assign n18990 = n18988 | n18989 ;
  assign n18991 = n12736 | n18990 ;
  assign n29156 = ~n18991 ;
  assign n18992 = x[11] & n29156 ;
  assign n18993 = n27892 & n18991 ;
  assign n18994 = n18992 | n18993 ;
  assign n18995 = n18987 & n18994 ;
  assign n19499 = n18987 | n18994 ;
  assign n29157 = ~n18995 ;
  assign n19500 = n29157 & n19499 ;
  assign n20061 = n19025 | n19027 ;
  assign n29158 = ~n19028 ;
  assign n20062 = n29158 & n20061 ;
  assign n20063 = n19485 & n20062 ;
  assign n20064 = n19028 | n20063 ;
  assign n20065 = n19009 | n19016 ;
  assign n20066 = n20064 & n20065 ;
  assign n20067 = n19018 | n20066 ;
  assign n20069 = n20067 & n20068 ;
  assign n20071 = n19005 | n20069 ;
  assign n29159 = ~n20071 ;
  assign n20072 = n19500 & n29159 ;
  assign n29160 = ~n19500 ;
  assign n20272 = n29160 & n20071 ;
  assign n20273 = n20072 | n20272 ;
  assign n29161 = ~n20271 ;
  assign n20842 = n29161 & n20273 ;
  assign n29162 = ~n20273 ;
  assign n21251 = n20271 & n29162 ;
  assign n21252 = n20842 | n21251 ;
  assign n21253 = n21250 | n21252 ;
  assign n21254 = n21250 & n21252 ;
  assign n29163 = ~n21254 ;
  assign n21427 = n21253 & n29163 ;
  assign n18416 = n2466 & n18392 ;
  assign n18333 = x[98] & n18329 ;
  assign n18555 = x[99] & n18514 ;
  assign n21428 = n18333 | n18555 ;
  assign n21429 = x[100] & n18327 ;
  assign n21430 = n21428 | n21429 ;
  assign n21431 = n18416 | n21430 ;
  assign n29164 = ~n21431 ;
  assign n21432 = x[5] & n29164 ;
  assign n21433 = n27813 & n21431 ;
  assign n21434 = n21432 | n21433 ;
  assign n21435 = n21427 & n21434 ;
  assign n21962 = n21427 | n21434 ;
  assign n29165 = ~n21435 ;
  assign n22252 = n29165 & n21962 ;
  assign n29166 = ~n21961 ;
  assign n22254 = n29166 & n22252 ;
  assign n29167 = ~n22252 ;
  assign n22444 = n21961 & n29167 ;
  assign n22445 = n22254 | n22444 ;
  assign n29168 = ~n22443 ;
  assign n22446 = n29168 & n22445 ;
  assign n29169 = ~n22445 ;
  assign n22448 = n22443 & n29169 ;
  assign n22449 = n22446 | n22448 ;
  assign n23003 = n22459 | n23002 ;
  assign n23004 = n22449 | n23003 ;
  assign n23005 = n22449 & n23003 ;
  assign n29170 = ~n23005 ;
  assign n168 = n23004 & n29170 ;
  assign n22447 = n22443 & n22445 ;
  assign n23006 = n22447 | n23005 ;
  assign n21963 = n21961 & n21962 ;
  assign n21964 = n21435 | n21963 ;
  assign n18435 = n2977 & n18392 ;
  assign n18384 = x[99] & n18329 ;
  assign n18550 = x[100] & n18514 ;
  assign n21417 = n18384 | n18550 ;
  assign n21418 = x[101] & n18327 ;
  assign n21419 = n21417 | n21418 ;
  assign n21420 = n18435 | n21419 ;
  assign n29171 = ~n21420 ;
  assign n21421 = x[5] & n29171 ;
  assign n21422 = n27813 & n21420 ;
  assign n21423 = n21421 | n21422 ;
  assign n20274 = n20271 & n20273 ;
  assign n21255 = n20274 | n21254 ;
  assign n15338 = n2841 & n15308 ;
  assign n15283 = x[96] & n15246 ;
  assign n17276 = x[97] & n16288 ;
  assign n20255 = n15283 | n17276 ;
  assign n20256 = x[98] & n15244 ;
  assign n20257 = n20255 | n20256 ;
  assign n20258 = n15338 | n20257 ;
  assign n29172 = ~n20258 ;
  assign n20259 = x[8] & n29172 ;
  assign n20260 = n27845 & n20258 ;
  assign n20261 = n20259 | n20260 ;
  assign n19497 = n19495 & n19496 ;
  assign n19498 = n19005 | n19497 ;
  assign n19501 = n19498 & n19500 ;
  assign n19502 = n18995 | n19501 ;
  assign n10564 = n1841 & n10542 ;
  assign n10496 = x[90] & n10481 ;
  assign n11909 = x[91] & n11232 ;
  assign n17728 = n10496 | n11909 ;
  assign n17729 = x[92] & n10479 ;
  assign n17730 = n17728 | n17729 ;
  assign n17731 = n10564 | n17730 ;
  assign n29173 = ~n17731 ;
  assign n17732 = x[14] & n29173 ;
  assign n17733 = n27956 & n17731 ;
  assign n17734 = n17732 | n17733 ;
  assign n17126 = n17123 & n17124 ;
  assign n17127 = n16788 | n17126 ;
  assign n7174 = n1213 & n7162 ;
  assign n7111 = x[84] & n7100 ;
  assign n7726 = x[85] & n7647 ;
  assign n15850 = n7111 | n7726 ;
  assign n15851 = x[86] & n7098 ;
  assign n15852 = n15850 | n15851 ;
  assign n15853 = n7174 | n15852 ;
  assign n29174 = ~n15853 ;
  assign n15854 = x[20] & n29174 ;
  assign n15855 = n28114 & n15853 ;
  assign n15856 = n15854 | n15855 ;
  assign n1273 = n452 & n1270 ;
  assign n341 = x[78] & n330 ;
  assign n441 = x[79] & n390 ;
  assign n13936 = n341 | n441 ;
  assign n13937 = x[80] & n322 ;
  assign n13938 = n13936 | n13937 ;
  assign n13939 = n1273 | n13938 ;
  assign n29175 = ~n13939 ;
  assign n13940 = x[26] & n29175 ;
  assign n13941 = n28342 & n13939 ;
  assign n13942 = n13940 | n13941 ;
  assign n13219 = n13210 & n13217 ;
  assign n13378 = n13219 | n13377 ;
  assign n12346 = n12337 & n12344 ;
  assign n12456 = n12346 | n12455 ;
  assign n4794 = n4041 & n4790 ;
  assign n3919 = x[69] & n3910 ;
  assign n4012 = x[70] & n3975 ;
  assign n11543 = n3919 | n4012 ;
  assign n11544 = x[71] & n3906 ;
  assign n11545 = n11543 | n11544 ;
  assign n11546 = n4794 | n11545 ;
  assign n29176 = ~n11546 ;
  assign n11547 = x[35] & n29176 ;
  assign n11548 = n28822 & n11546 ;
  assign n11549 = n11547 | n11548 ;
  assign n11023 = n11014 & n11021 ;
  assign n11024 = n11012 | n11023 ;
  assign n6412 = n3574 & n6408 ;
  assign n3462 = x[66] & n3443 ;
  assign n3520 = x[67] & n3508 ;
  assign n10982 = n3462 | n3520 ;
  assign n10983 = x[68] & n3439 ;
  assign n10984 = n10982 | n10983 ;
  assign n10985 = n6412 | n10984 ;
  assign n10986 = x[38] | n10985 ;
  assign n10987 = x[38] & n10985 ;
  assign n29177 = ~n10987 ;
  assign n10988 = n10986 & n29177 ;
  assign n29178 = ~n10239 ;
  assign n10240 = x[41] & n29178 ;
  assign n27723 = x[40] & x[41] ;
  assign n3025 = x[40] | x[41] ;
  assign n29179 = ~n27723 ;
  assign n3026 = n29179 & n3025 ;
  assign n3162 = n3024 & n3026 ;
  assign n6441 = n3162 & n6437 ;
  assign n29180 = ~n3026 ;
  assign n3027 = n3024 & n29180 ;
  assign n10241 = x[65] & n3027 ;
  assign n27725 = x[39] & x[40] ;
  assign n3028 = x[39] | x[40] ;
  assign n29181 = ~n27725 ;
  assign n3029 = n29181 & n3028 ;
  assign n29182 = ~n3024 ;
  assign n3096 = n29182 & n3029 ;
  assign n10242 = x[64] & n3096 ;
  assign n10243 = n10241 | n10242 ;
  assign n10244 = n6441 | n10243 ;
  assign n29183 = ~n10244 ;
  assign n10245 = x[41] & n29183 ;
  assign n29184 = ~x[41] ;
  assign n10246 = n29184 & n10244 ;
  assign n10247 = n10245 | n10246 ;
  assign n29185 = ~n10247 ;
  assign n10248 = n10240 & n29185 ;
  assign n29186 = ~n10240 ;
  assign n10989 = n29186 & n10247 ;
  assign n10990 = n10248 | n10989 ;
  assign n10991 = n10988 & n10990 ;
  assign n11025 = n10988 | n10990 ;
  assign n29187 = ~n10991 ;
  assign n11026 = n29187 & n11025 ;
  assign n29188 = ~n11024 ;
  assign n11027 = n29188 & n11026 ;
  assign n29189 = ~n11026 ;
  assign n11550 = n11024 & n29189 ;
  assign n11551 = n11027 | n11550 ;
  assign n29190 = ~n11549 ;
  assign n11552 = n29190 & n11551 ;
  assign n29191 = ~n11551 ;
  assign n11554 = n11549 & n29191 ;
  assign n11555 = n11552 | n11554 ;
  assign n11633 = n11567 & n11631 ;
  assign n11634 = n11565 | n11633 ;
  assign n29192 = ~n11634 ;
  assign n11635 = n11555 & n29192 ;
  assign n29193 = ~n11555 ;
  assign n12326 = n29193 & n11634 ;
  assign n12327 = n11635 | n12326 ;
  assign n2724 = n779 & n2722 ;
  assign n677 = x[72] & n663 ;
  assign n768 = x[73] & n720 ;
  assign n12328 = n677 | n768 ;
  assign n12329 = x[74] & n652 ;
  assign n12330 = n12328 | n12329 ;
  assign n12331 = n2724 | n12330 ;
  assign n29194 = ~n12331 ;
  assign n12332 = x[32] & n29194 ;
  assign n12333 = n28658 & n12331 ;
  assign n12334 = n12332 | n12333 ;
  assign n12335 = n12327 & n12334 ;
  assign n12457 = n12327 | n12334 ;
  assign n29195 = ~n12335 ;
  assign n13197 = n29195 & n12457 ;
  assign n29196 = ~n13197 ;
  assign n13198 = n12456 & n29196 ;
  assign n12458 = n12456 & n12457 ;
  assign n12459 = n12335 | n12458 ;
  assign n29197 = ~n12459 ;
  assign n13199 = n12457 & n29197 ;
  assign n13200 = n13198 | n13199 ;
  assign n4660 = n1775 & n4632 ;
  assign n4546 = x[75] & n4514 ;
  assign n4594 = x[76] & n4572 ;
  assign n13201 = n4546 | n4594 ;
  assign n13202 = x[77] & n4504 ;
  assign n13203 = n13201 | n13202 ;
  assign n13204 = n4660 | n13203 ;
  assign n29198 = ~n13204 ;
  assign n13205 = x[29] & n29198 ;
  assign n13206 = n28483 & n13204 ;
  assign n13207 = n13205 | n13206 ;
  assign n29199 = ~n13207 ;
  assign n13208 = n13200 & n29199 ;
  assign n29200 = ~n13200 ;
  assign n13379 = n29200 & n13207 ;
  assign n13380 = n13208 | n13379 ;
  assign n13381 = n13378 & n13380 ;
  assign n13943 = n13378 | n13380 ;
  assign n29201 = ~n13381 ;
  assign n13944 = n29201 & n13943 ;
  assign n29202 = ~n13942 ;
  assign n13946 = n29202 & n13944 ;
  assign n29203 = ~n13944 ;
  assign n13947 = n13942 & n29203 ;
  assign n13948 = n13946 | n13947 ;
  assign n29204 = ~n13374 ;
  assign n13375 = n13221 & n29204 ;
  assign n29205 = ~n13221 ;
  assign n13956 = n29205 & n13374 ;
  assign n13957 = n13375 | n13956 ;
  assign n13958 = n13955 & n13957 ;
  assign n14161 = n13967 & n14160 ;
  assign n14162 = n13968 | n14161 ;
  assign n14164 = n13955 & n14163 ;
  assign n14166 = n13955 | n14163 ;
  assign n29206 = ~n14164 ;
  assign n14167 = n29206 & n14166 ;
  assign n14168 = n14162 & n14167 ;
  assign n14169 = n13958 | n14168 ;
  assign n14170 = n13948 | n14169 ;
  assign n14171 = n13948 & n14169 ;
  assign n29207 = ~n14171 ;
  assign n14840 = n14170 & n29207 ;
  assign n5312 = n1057 & n5302 ;
  assign n5269 = x[81] & n5240 ;
  assign n6255 = x[82] & n6179 ;
  assign n14841 = n5269 | n6255 ;
  assign n14842 = x[83] & n5238 ;
  assign n14843 = n14841 | n14842 ;
  assign n14844 = n5312 | n14843 ;
  assign n29208 = ~n14844 ;
  assign n14845 = x[23] & n29208 ;
  assign n14846 = n28221 & n14844 ;
  assign n14847 = n14845 | n14846 ;
  assign n29209 = ~n14847 ;
  assign n14848 = n14840 & n29209 ;
  assign n29210 = ~n14840 ;
  assign n15732 = n29210 & n14847 ;
  assign n15733 = n14848 | n15732 ;
  assign n15786 = n14864 | n15785 ;
  assign n15788 = n15733 | n15786 ;
  assign n15789 = n15733 & n15786 ;
  assign n29211 = ~n15789 ;
  assign n15859 = n15788 & n29211 ;
  assign n29212 = ~n15856 ;
  assign n15860 = n29212 & n15859 ;
  assign n29213 = ~n15859 ;
  assign n15861 = n15856 & n29213 ;
  assign n15862 = n15860 | n15861 ;
  assign n16164 = n15886 | n16163 ;
  assign n16165 = n15875 & n16164 ;
  assign n16166 = n15873 | n16165 ;
  assign n16167 = n15862 | n16166 ;
  assign n16168 = n15862 & n16166 ;
  assign n29214 = ~n16168 ;
  assign n16763 = n16167 & n29214 ;
  assign n8721 = n1453 & n8706 ;
  assign n8660 = x[87] & n8645 ;
  assign n9881 = x[88] & n9278 ;
  assign n16764 = n8660 | n9881 ;
  assign n16765 = x[89] & n8643 ;
  assign n16766 = n16764 | n16765 ;
  assign n16767 = n8721 | n16766 ;
  assign n29215 = ~n16767 ;
  assign n16768 = x[17] & n29215 ;
  assign n16769 = n28039 & n16767 ;
  assign n16770 = n16768 | n16769 ;
  assign n29216 = ~n16770 ;
  assign n16771 = n16763 & n29216 ;
  assign n29217 = ~n16763 ;
  assign n17454 = n29217 & n16770 ;
  assign n17455 = n16771 | n17454 ;
  assign n17457 = n17127 | n17455 ;
  assign n17458 = n17127 & n17455 ;
  assign n29218 = ~n17458 ;
  assign n18206 = n17457 & n29218 ;
  assign n29219 = ~n17734 ;
  assign n18207 = n29219 & n18206 ;
  assign n29220 = ~n18206 ;
  assign n18209 = n17734 & n29220 ;
  assign n18210 = n18207 | n18209 ;
  assign n17747 = n17744 & n17746 ;
  assign n18724 = n17747 | n18723 ;
  assign n29221 = ~n18210 ;
  assign n18725 = n29221 & n18724 ;
  assign n29222 = ~n18724 ;
  assign n18977 = n18210 & n29222 ;
  assign n18978 = n18725 | n18977 ;
  assign n12733 = n2152 & n12695 ;
  assign n12639 = x[93] & n12633 ;
  assign n14372 = x[94] & n13533 ;
  assign n18979 = n12639 | n14372 ;
  assign n18980 = x[95] & n12631 ;
  assign n18981 = n18979 | n18980 ;
  assign n18982 = n12733 | n18981 ;
  assign n29223 = ~n18982 ;
  assign n18983 = x[11] & n29223 ;
  assign n18984 = n27892 & n18982 ;
  assign n18985 = n18983 | n18984 ;
  assign n18986 = n18978 & n18985 ;
  assign n19503 = n18978 | n18985 ;
  assign n29224 = ~n18986 ;
  assign n20075 = n29224 & n19503 ;
  assign n29225 = ~n19502 ;
  assign n20077 = n29225 & n20075 ;
  assign n29226 = ~n20075 ;
  assign n20262 = n19502 & n29226 ;
  assign n20263 = n20077 | n20262 ;
  assign n20264 = n20261 & n20263 ;
  assign n20847 = n20261 | n20263 ;
  assign n29227 = ~n20264 ;
  assign n21256 = n29227 & n20847 ;
  assign n21257 = n21255 & n21256 ;
  assign n21965 = n21255 | n21256 ;
  assign n29228 = ~n21257 ;
  assign n21966 = n29228 & n21965 ;
  assign n29229 = ~n21423 ;
  assign n21968 = n29229 & n21966 ;
  assign n29230 = ~n21966 ;
  assign n22256 = n21423 & n29230 ;
  assign n22257 = n21968 | n22256 ;
  assign n29231 = ~n22257 ;
  assign n22258 = n21964 & n29231 ;
  assign n29232 = ~n21964 ;
  assign n22426 = n29232 & n22257 ;
  assign n22427 = n22258 | n22426 ;
  assign n573 = n571 & n572 ;
  assign n574 = n27624 | n573 ;
  assign n25228 = x[103] & x[104] ;
  assign n575 = x[103] | x[104] ;
  assign n29233 = ~n25228 ;
  assign n2998 = n29233 & n575 ;
  assign n2999 = n574 & n2998 ;
  assign n3000 = n574 | n2998 ;
  assign n29234 = ~n2999 ;
  assign n3001 = n29234 & n3000 ;
  assign n19716 = n3001 & n19656 ;
  assign n19782 = x[102] & n19723 ;
  assign n19884 = x[103] & n19829 ;
  assign n22428 = n19782 | n19884 ;
  assign n22429 = x[104] & n19655 ;
  assign n22430 = n22428 | n22429 ;
  assign n22431 = n19716 | n22430 ;
  assign n29235 = ~n22431 ;
  assign n22432 = x[2] & n29235 ;
  assign n22433 = n27790 & n22431 ;
  assign n22434 = n22432 | n22433 ;
  assign n22435 = n22427 | n22434 ;
  assign n22436 = n22427 & n22434 ;
  assign n29236 = ~n22436 ;
  assign n23007 = n22435 & n29236 ;
  assign n23008 = n23006 & n23007 ;
  assign n27681 = n23006 | n23007 ;
  assign n29237 = ~n23008 ;
  assign n169 = n29237 & n27681 ;
  assign n23009 = n22436 | n23008 ;
  assign n20840 = n20838 & n20839 ;
  assign n20841 = n20284 | n20840 ;
  assign n20843 = n20271 | n20273 ;
  assign n29238 = ~n20274 ;
  assign n20844 = n29238 & n20843 ;
  assign n20845 = n20841 & n20844 ;
  assign n20846 = n20274 | n20845 ;
  assign n29239 = ~n20846 ;
  assign n21258 = n29239 & n21256 ;
  assign n29240 = ~n21256 ;
  assign n21424 = n20846 & n29240 ;
  assign n21425 = n21258 | n21424 ;
  assign n21426 = n21423 & n21425 ;
  assign n21967 = n21423 & n21966 ;
  assign n21969 = n21423 | n21966 ;
  assign n29241 = ~n21967 ;
  assign n21970 = n29241 & n21969 ;
  assign n21971 = n21964 & n21970 ;
  assign n21972 = n21426 | n21971 ;
  assign n20848 = n20846 & n20847 ;
  assign n20849 = n20264 | n20848 ;
  assign n15324 = n2313 & n15308 ;
  assign n15300 = x[97] & n15246 ;
  assign n17293 = x[98] & n16288 ;
  assign n20245 = n15300 | n17293 ;
  assign n20246 = x[99] & n15244 ;
  assign n20247 = n20245 | n20246 ;
  assign n20248 = n15324 | n20247 ;
  assign n29242 = ~n20248 ;
  assign n20249 = x[8] & n29242 ;
  assign n20250 = n27845 & n20248 ;
  assign n20251 = n20249 | n20250 ;
  assign n12754 = n2000 & n12695 ;
  assign n12657 = x[94] & n12633 ;
  assign n14362 = x[95] & n13533 ;
  assign n18967 = n12657 | n14362 ;
  assign n18968 = x[96] & n12631 ;
  assign n18969 = n18967 | n18968 ;
  assign n18970 = n12754 | n18969 ;
  assign n29243 = ~n18970 ;
  assign n18971 = x[11] & n29243 ;
  assign n18972 = n27892 & n18970 ;
  assign n18973 = n18971 | n18972 ;
  assign n13945 = n13942 & n13944 ;
  assign n14698 = n13942 | n13944 ;
  assign n29244 = ~n13945 ;
  assign n14699 = n29244 & n14698 ;
  assign n29245 = ~n14169 ;
  assign n14700 = n29245 & n14699 ;
  assign n29246 = ~n14699 ;
  assign n14850 = n14169 & n29246 ;
  assign n14851 = n14700 | n14850 ;
  assign n14852 = n14847 | n14851 ;
  assign n14853 = n14847 & n14851 ;
  assign n29247 = ~n14853 ;
  assign n14854 = n14852 & n29247 ;
  assign n29248 = ~n15786 ;
  assign n15787 = n14854 & n29248 ;
  assign n29249 = ~n14854 ;
  assign n15848 = n29249 & n15786 ;
  assign n15849 = n15787 | n15848 ;
  assign n15857 = n15849 | n15856 ;
  assign n15858 = n15849 & n15856 ;
  assign n29250 = ~n15858 ;
  assign n16409 = n15857 & n29250 ;
  assign n29251 = ~n16166 ;
  assign n16410 = n29251 & n16409 ;
  assign n29252 = ~n16409 ;
  assign n16773 = n16166 & n29252 ;
  assign n16774 = n16410 | n16773 ;
  assign n16775 = n16770 | n16774 ;
  assign n16776 = n16770 & n16774 ;
  assign n29253 = ~n16776 ;
  assign n16777 = n16775 & n29253 ;
  assign n29254 = ~n17127 ;
  assign n17456 = n16777 & n29254 ;
  assign n29255 = ~n16777 ;
  assign n17735 = n29255 & n17127 ;
  assign n17736 = n17456 | n17735 ;
  assign n17737 = n17734 & n17736 ;
  assign n18198 = n17825 | n17832 ;
  assign n18199 = n18197 & n18198 ;
  assign n18200 = n17834 | n18199 ;
  assign n18202 = n17744 | n17746 ;
  assign n29256 = ~n17747 ;
  assign n18203 = n29256 & n18202 ;
  assign n18204 = n18200 & n18203 ;
  assign n18205 = n17747 | n18204 ;
  assign n18211 = n18205 & n18210 ;
  assign n18212 = n17737 | n18211 ;
  assign n10565 = n1685 & n10542 ;
  assign n10492 = x[91] & n10481 ;
  assign n11878 = x[92] & n11232 ;
  assign n17718 = n10492 | n11878 ;
  assign n17719 = x[93] & n10479 ;
  assign n17720 = n17718 | n17719 ;
  assign n17721 = n10565 | n17720 ;
  assign n29257 = ~n17721 ;
  assign n17722 = x[14] & n29257 ;
  assign n17723 = n27956 & n17721 ;
  assign n17724 = n17722 | n17723 ;
  assign n17459 = n16776 | n17458 ;
  assign n16169 = n15858 | n16168 ;
  assign n5348 = n1293 & n5302 ;
  assign n5273 = x[82] & n5240 ;
  assign n6232 = x[83] & n6179 ;
  assign n14827 = n5273 | n6232 ;
  assign n14828 = x[84] & n5238 ;
  assign n14829 = n14827 | n14828 ;
  assign n14830 = n5348 | n14829 ;
  assign n29258 = ~n14830 ;
  assign n14831 = x[23] & n29258 ;
  assign n14832 = n28221 & n14830 ;
  assign n14833 = n14831 | n14832 ;
  assign n14172 = n13945 | n14171 ;
  assign n1030 = n452 & n1029 ;
  assign n342 = x[79] & n330 ;
  assign n433 = x[80] & n390 ;
  assign n13926 = n342 | n433 ;
  assign n13927 = x[81] & n322 ;
  assign n13928 = n13926 | n13927 ;
  assign n13929 = n1030 | n13928 ;
  assign n29259 = ~n13929 ;
  assign n13930 = x[26] & n29259 ;
  assign n13931 = n28342 & n13929 ;
  assign n13932 = n13930 | n13931 ;
  assign n13209 = n13200 & n13207 ;
  assign n13382 = n13209 | n13381 ;
  assign n4637 = n2084 & n4632 ;
  assign n4562 = x[76] & n4514 ;
  assign n4578 = x[77] & n4572 ;
  assign n13187 = n4562 | n4578 ;
  assign n13188 = x[78] & n4504 ;
  assign n13189 = n13187 | n13188 ;
  assign n13190 = n4637 | n13189 ;
  assign n29260 = ~n13190 ;
  assign n13191 = x[29] & n29260 ;
  assign n13192 = n28483 & n13190 ;
  assign n13193 = n13191 | n13192 ;
  assign n11553 = n11549 & n11551 ;
  assign n11636 = n11555 & n11634 ;
  assign n11637 = n11553 | n11636 ;
  assign n4054 = n3701 & n4041 ;
  assign n3947 = x[70] & n3910 ;
  assign n3985 = x[71] & n3975 ;
  assign n11532 = n3947 | n3985 ;
  assign n11533 = x[72] & n3906 ;
  assign n11534 = n11532 | n11533 ;
  assign n11535 = n4054 | n11534 ;
  assign n29261 = ~n11535 ;
  assign n11536 = x[35] & n29261 ;
  assign n11537 = n28822 & n11535 ;
  assign n11538 = n11536 | n11537 ;
  assign n11028 = n11024 & n11026 ;
  assign n11029 = n10991 | n11028 ;
  assign n10249 = n10240 & n10247 ;
  assign n6473 = n3162 & n6466 ;
  assign n3030 = n29182 & n3026 ;
  assign n29262 = ~n3029 ;
  assign n3031 = n29262 & n3030 ;
  assign n3040 = x[64] & n3031 ;
  assign n3101 = x[65] & n3096 ;
  assign n10250 = n3040 | n3101 ;
  assign n10251 = x[66] & n3027 ;
  assign n10252 = n10250 | n10251 ;
  assign n10253 = n6473 | n10252 ;
  assign n29263 = ~n10253 ;
  assign n10254 = x[41] & n29263 ;
  assign n10255 = n29184 & n10253 ;
  assign n10256 = n10254 | n10255 ;
  assign n29264 = ~n10256 ;
  assign n10257 = n10249 & n29264 ;
  assign n29265 = ~n10249 ;
  assign n10971 = n29265 & n10256 ;
  assign n10972 = n10257 | n10971 ;
  assign n6381 = n3574 & n6379 ;
  assign n3451 = x[67] & n3443 ;
  assign n3516 = x[68] & n3508 ;
  assign n10973 = n3451 | n3516 ;
  assign n10974 = x[69] & n3439 ;
  assign n10975 = n10973 | n10974 ;
  assign n10976 = n6381 | n10975 ;
  assign n29266 = ~n10976 ;
  assign n10977 = x[38] & n29266 ;
  assign n10978 = n28996 & n10976 ;
  assign n10979 = n10977 | n10978 ;
  assign n29267 = ~n10979 ;
  assign n10980 = n10972 & n29267 ;
  assign n29268 = ~n10972 ;
  assign n11030 = n29268 & n10979 ;
  assign n11031 = n10980 | n11030 ;
  assign n29269 = ~n11031 ;
  assign n11032 = n11029 & n29269 ;
  assign n29270 = ~n11029 ;
  assign n11539 = n29270 & n11031 ;
  assign n11540 = n11032 | n11539 ;
  assign n29271 = ~n11538 ;
  assign n11541 = n29271 & n11540 ;
  assign n29272 = ~n11540 ;
  assign n11638 = n11538 & n29272 ;
  assign n11639 = n11541 | n11638 ;
  assign n29273 = ~n11639 ;
  assign n11640 = n11637 & n29273 ;
  assign n29274 = ~n11637 ;
  assign n12315 = n29274 & n11639 ;
  assign n12316 = n11640 | n12315 ;
  assign n3293 = n779 & n3289 ;
  assign n701 = x[73] & n663 ;
  assign n767 = x[74] & n720 ;
  assign n12317 = n701 | n767 ;
  assign n12318 = x[75] & n652 ;
  assign n12319 = n12317 | n12318 ;
  assign n12320 = n3293 | n12319 ;
  assign n29275 = ~n12320 ;
  assign n12321 = x[32] & n29275 ;
  assign n12322 = n28658 & n12320 ;
  assign n12323 = n12321 | n12322 ;
  assign n12324 = n12316 | n12323 ;
  assign n12325 = n12316 & n12323 ;
  assign n29276 = ~n12325 ;
  assign n12460 = n12324 & n29276 ;
  assign n12461 = n29197 & n12460 ;
  assign n29277 = ~n12460 ;
  assign n13194 = n12459 & n29277 ;
  assign n13195 = n12461 | n13194 ;
  assign n13196 = n13193 & n13195 ;
  assign n13383 = n13193 | n13195 ;
  assign n29278 = ~n13196 ;
  assign n13781 = n29278 & n13383 ;
  assign n29279 = ~n13382 ;
  assign n13783 = n29279 & n13781 ;
  assign n29280 = ~n13781 ;
  assign n13933 = n13382 & n29280 ;
  assign n13934 = n13783 | n13933 ;
  assign n13935 = n13932 & n13934 ;
  assign n14173 = n13932 | n13934 ;
  assign n29281 = ~n13935 ;
  assign n14174 = n29281 & n14173 ;
  assign n14175 = n14172 & n14174 ;
  assign n14834 = n14172 | n14174 ;
  assign n29282 = ~n14175 ;
  assign n14835 = n29282 & n14834 ;
  assign n29283 = ~n14833 ;
  assign n14837 = n29283 & n14835 ;
  assign n29284 = ~n14835 ;
  assign n14838 = n14833 & n29284 ;
  assign n14839 = n14837 | n14838 ;
  assign n14849 = n14840 & n14847 ;
  assign n15102 = n14887 | n15101 ;
  assign n15103 = n14877 & n15102 ;
  assign n15104 = n14874 | n15103 ;
  assign n15105 = n14863 & n15104 ;
  assign n15106 = n14864 | n15105 ;
  assign n15107 = n14854 & n15106 ;
  assign n15108 = n14849 | n15107 ;
  assign n15109 = n14839 | n15108 ;
  assign n15110 = n14839 & n15108 ;
  assign n29285 = ~n15110 ;
  assign n15839 = n15109 & n29285 ;
  assign n7175 = n1522 & n7162 ;
  assign n7112 = x[85] & n7100 ;
  assign n7686 = x[86] & n7647 ;
  assign n15840 = n7112 | n7686 ;
  assign n15841 = x[87] & n7098 ;
  assign n15842 = n15840 | n15841 ;
  assign n15843 = n7175 | n15842 ;
  assign n29286 = ~n15843 ;
  assign n15844 = x[20] & n29286 ;
  assign n15845 = n28114 & n15843 ;
  assign n15846 = n15844 | n15845 ;
  assign n15847 = n15839 & n15846 ;
  assign n14836 = n14833 & n14835 ;
  assign n15729 = n14833 | n14835 ;
  assign n29287 = ~n14836 ;
  assign n15730 = n29287 & n15729 ;
  assign n29288 = ~n15108 ;
  assign n15731 = n29288 & n15730 ;
  assign n29289 = ~n15730 ;
  assign n16405 = n15108 & n29289 ;
  assign n16406 = n15731 | n16405 ;
  assign n16473 = n15846 | n16406 ;
  assign n29290 = ~n15847 ;
  assign n16750 = n29290 & n16473 ;
  assign n29291 = ~n16750 ;
  assign n16751 = n16169 & n29291 ;
  assign n16407 = n15846 & n16406 ;
  assign n16408 = n15856 & n15859 ;
  assign n29292 = ~n15871 ;
  assign n15872 = n15864 & n29292 ;
  assign n29293 = ~n15864 ;
  assign n16411 = n29293 & n15871 ;
  assign n16412 = n15872 | n16411 ;
  assign n16469 = n16412 & n16467 ;
  assign n16470 = n15873 | n16469 ;
  assign n16471 = n16409 & n16470 ;
  assign n16472 = n16408 | n16471 ;
  assign n16474 = n16472 & n16473 ;
  assign n16475 = n16407 | n16474 ;
  assign n29294 = ~n16475 ;
  assign n16752 = n16473 & n29294 ;
  assign n16753 = n16751 | n16752 ;
  assign n8756 = n1482 & n8706 ;
  assign n8664 = x[88] & n8645 ;
  assign n9878 = x[89] & n9278 ;
  assign n16754 = n8664 | n9878 ;
  assign n16755 = x[90] & n8643 ;
  assign n16756 = n16754 | n16755 ;
  assign n16757 = n8756 | n16756 ;
  assign n29295 = ~n16757 ;
  assign n16758 = x[17] & n29295 ;
  assign n16759 = n28039 & n16757 ;
  assign n16760 = n16758 | n16759 ;
  assign n29296 = ~n16760 ;
  assign n16761 = n16753 & n29296 ;
  assign n29297 = ~n16753 ;
  assign n17460 = n29297 & n16760 ;
  assign n17461 = n16761 | n17460 ;
  assign n17462 = n17459 & n17461 ;
  assign n17725 = n17459 | n17461 ;
  assign n29298 = ~n17462 ;
  assign n17726 = n29298 & n17725 ;
  assign n17727 = n17724 & n17726 ;
  assign n18213 = n17724 | n17726 ;
  assign n29299 = ~n17727 ;
  assign n18214 = n29299 & n18213 ;
  assign n18215 = n18212 & n18214 ;
  assign n18974 = n18212 | n18214 ;
  assign n29300 = ~n18215 ;
  assign n18975 = n29300 & n18974 ;
  assign n18976 = n18973 & n18975 ;
  assign n19506 = n18973 | n18975 ;
  assign n29301 = ~n18976 ;
  assign n19507 = n29301 & n19506 ;
  assign n20073 = n19499 & n20071 ;
  assign n20074 = n18995 | n20073 ;
  assign n20076 = n20074 & n20075 ;
  assign n20078 = n18986 | n20076 ;
  assign n29302 = ~n20078 ;
  assign n20079 = n19507 & n29302 ;
  assign n29303 = ~n19507 ;
  assign n20252 = n29303 & n20078 ;
  assign n20253 = n20079 | n20252 ;
  assign n29304 = ~n20251 ;
  assign n20850 = n29304 & n20253 ;
  assign n29305 = ~n20253 ;
  assign n21260 = n20251 & n29305 ;
  assign n21261 = n20850 | n21260 ;
  assign n29306 = ~n21261 ;
  assign n21262 = n20849 & n29306 ;
  assign n29307 = ~n20849 ;
  assign n21407 = n29307 & n21261 ;
  assign n21408 = n21262 | n21407 ;
  assign n18446 = n2867 & n18392 ;
  assign n18381 = x[100] & n18329 ;
  assign n18561 = x[101] & n18514 ;
  assign n21409 = n18381 | n18561 ;
  assign n21410 = x[102] & n18327 ;
  assign n21411 = n21409 | n21410 ;
  assign n21412 = n18446 | n21411 ;
  assign n29308 = ~n21412 ;
  assign n21413 = x[5] & n29308 ;
  assign n21414 = n27813 & n21412 ;
  assign n21415 = n21413 | n21414 ;
  assign n21416 = n21408 & n21415 ;
  assign n21259 = n20264 | n21257 ;
  assign n21263 = n21259 | n21261 ;
  assign n21264 = n21259 & n21261 ;
  assign n29309 = ~n21264 ;
  assign n21973 = n21263 & n29309 ;
  assign n21974 = n21415 | n21973 ;
  assign n29310 = ~n21416 ;
  assign n22261 = n29310 & n21974 ;
  assign n29311 = ~n21972 ;
  assign n22263 = n29311 & n22261 ;
  assign n29312 = ~n22261 ;
  assign n22415 = n21972 & n29312 ;
  assign n22416 = n22263 | n22415 ;
  assign n576 = n574 & n575 ;
  assign n577 = n25228 | n576 ;
  assign n27622 = x[104] & x[105] ;
  assign n578 = x[104] | x[105] ;
  assign n29313 = ~n27622 ;
  assign n3406 = n29313 & n578 ;
  assign n3407 = n577 | n3406 ;
  assign n3408 = n577 & n3406 ;
  assign n29314 = ~n3408 ;
  assign n3409 = n3407 & n29314 ;
  assign n19682 = n3409 & n19656 ;
  assign n19781 = x[103] & n19723 ;
  assign n19855 = x[104] & n19829 ;
  assign n22417 = n19781 | n19855 ;
  assign n22418 = x[105] & n19655 ;
  assign n22419 = n22417 | n22418 ;
  assign n22420 = n19682 | n22419 ;
  assign n29315 = ~n22420 ;
  assign n22421 = x[2] & n29315 ;
  assign n22422 = n27790 & n22420 ;
  assign n22423 = n22421 | n22422 ;
  assign n22424 = n22416 | n22423 ;
  assign n22425 = n22416 & n22423 ;
  assign n29316 = ~n22425 ;
  assign n23010 = n22424 & n29316 ;
  assign n23011 = n23009 | n23010 ;
  assign n23012 = n23009 & n23010 ;
  assign n29317 = ~n23012 ;
  assign n170 = n23011 & n29317 ;
  assign n22102 = n21415 & n21973 ;
  assign n22246 = n21952 & n22244 ;
  assign n22247 = n21468 | n22246 ;
  assign n22248 = n22104 & n22247 ;
  assign n22249 = n21455 | n22248 ;
  assign n22250 = n21958 & n22249 ;
  assign n22251 = n21445 | n22250 ;
  assign n22253 = n22251 & n22252 ;
  assign n22255 = n21435 | n22253 ;
  assign n22259 = n22255 & n22257 ;
  assign n22260 = n21426 | n22259 ;
  assign n22262 = n22260 & n22261 ;
  assign n22264 = n22102 | n22262 ;
  assign n18453 = n2626 & n18392 ;
  assign n18378 = x[101] & n18329 ;
  assign n18573 = x[102] & n18514 ;
  assign n21397 = n18378 | n18573 ;
  assign n21398 = x[103] & n18327 ;
  assign n21399 = n21397 | n21398 ;
  assign n21400 = n18453 | n21399 ;
  assign n29318 = ~n21400 ;
  assign n21401 = x[5] & n29318 ;
  assign n21402 = n27813 & n21400 ;
  assign n21403 = n21401 | n21402 ;
  assign n20254 = n20251 & n20253 ;
  assign n21265 = n20254 | n21264 ;
  assign n19504 = n19502 & n19503 ;
  assign n19505 = n18986 | n19504 ;
  assign n19508 = n19505 & n19507 ;
  assign n19509 = n18976 | n19508 ;
  assign n12729 = n2438 & n12695 ;
  assign n12687 = x[95] & n12633 ;
  assign n14404 = x[96] & n13533 ;
  assign n18957 = n12687 | n14404 ;
  assign n18958 = x[97] & n12631 ;
  assign n18959 = n18957 | n18958 ;
  assign n18960 = n12729 | n18959 ;
  assign n29319 = ~n18960 ;
  assign n18961 = x[11] & n29319 ;
  assign n18962 = n27892 & n18960 ;
  assign n18963 = n18961 | n18962 ;
  assign n18216 = n17727 | n18215 ;
  assign n16762 = n16753 & n16760 ;
  assign n17463 = n16762 | n17462 ;
  assign n8725 = n2046 & n8706 ;
  assign n8662 = x[89] & n8645 ;
  assign n9886 = x[90] & n9278 ;
  assign n16740 = n8662 | n9886 ;
  assign n16741 = x[91] & n8643 ;
  assign n16742 = n16740 | n16741 ;
  assign n16743 = n8725 | n16742 ;
  assign n29320 = ~n16743 ;
  assign n16744 = x[17] & n29320 ;
  assign n16745 = n28039 & n16743 ;
  assign n16746 = n16744 | n16745 ;
  assign n16170 = n15839 | n15846 ;
  assign n16171 = n16169 & n16170 ;
  assign n16172 = n15847 | n16171 ;
  assign n5332 = n1239 & n5302 ;
  assign n5252 = x[83] & n5240 ;
  assign n6233 = x[84] & n6179 ;
  assign n14814 = n5252 | n6233 ;
  assign n14815 = x[85] & n5238 ;
  assign n14816 = n14814 | n14815 ;
  assign n14817 = n5332 | n14816 ;
  assign n29321 = ~n14817 ;
  assign n14818 = x[23] & n29321 ;
  assign n14819 = n28221 & n14817 ;
  assign n14820 = n14818 | n14819 ;
  assign n14176 = n13935 | n14175 ;
  assign n13384 = n13382 & n13383 ;
  assign n13385 = n13196 | n13384 ;
  assign n12462 = n12459 & n12460 ;
  assign n12463 = n12325 | n12462 ;
  assign n2752 = n779 & n2750 ;
  assign n665 = x[74] & n663 ;
  assign n766 = x[75] & n720 ;
  assign n12305 = n665 | n766 ;
  assign n12306 = x[76] & n652 ;
  assign n12307 = n12305 | n12306 ;
  assign n12308 = n2752 | n12307 ;
  assign n29322 = ~n12308 ;
  assign n12309 = x[32] & n29322 ;
  assign n12310 = n28658 & n12308 ;
  assign n12311 = n12309 | n12310 ;
  assign n11542 = n11538 & n11540 ;
  assign n11641 = n11637 & n11639 ;
  assign n11642 = n11542 | n11641 ;
  assign n5980 = n3574 & n5976 ;
  assign n3455 = x[68] & n3443 ;
  assign n3518 = x[69] & n3508 ;
  assign n10959 = n3455 | n3518 ;
  assign n10960 = x[70] & n3439 ;
  assign n10961 = n10959 | n10960 ;
  assign n10962 = n5980 | n10961 ;
  assign n29323 = ~n10962 ;
  assign n10963 = x[38] & n29323 ;
  assign n10964 = n28996 & n10962 ;
  assign n10965 = n10963 | n10964 ;
  assign n27706 = x[41] & x[42] ;
  assign n2484 = x[41] | x[42] ;
  assign n29324 = ~n27706 ;
  assign n2485 = n29324 & n2484 ;
  assign n9557 = x[64] & n2485 ;
  assign n10258 = n10249 & n10256 ;
  assign n10259 = n9557 & n10258 ;
  assign n10260 = n9557 | n10258 ;
  assign n29325 = ~n10259 ;
  assign n10261 = n29325 & n10260 ;
  assign n6501 = n3162 & n6494 ;
  assign n3039 = x[65] & n3031 ;
  assign n3144 = x[66] & n3096 ;
  assign n10262 = n3039 | n3144 ;
  assign n10263 = x[67] & n3027 ;
  assign n10264 = n10262 | n10263 ;
  assign n10265 = n6501 | n10264 ;
  assign n29326 = ~n10265 ;
  assign n10266 = x[41] & n29326 ;
  assign n10267 = n29184 & n10265 ;
  assign n10268 = n10266 | n10267 ;
  assign n29327 = ~n10268 ;
  assign n10269 = n10261 & n29327 ;
  assign n29328 = ~n10261 ;
  assign n10966 = n29328 & n10268 ;
  assign n10967 = n10269 | n10966 ;
  assign n10968 = n10965 & n10967 ;
  assign n10969 = n10965 | n10967 ;
  assign n29329 = ~n10968 ;
  assign n10970 = n29329 & n10969 ;
  assign n10981 = n10972 & n10979 ;
  assign n11033 = n11029 & n11031 ;
  assign n11034 = n10981 | n11033 ;
  assign n29330 = ~n11034 ;
  assign n11035 = n10970 & n29330 ;
  assign n29331 = ~n10970 ;
  assign n11522 = n29331 & n11034 ;
  assign n11523 = n11035 | n11522 ;
  assign n4044 = n3733 & n4041 ;
  assign n3920 = x[71] & n3910 ;
  assign n4005 = x[72] & n3975 ;
  assign n11524 = n3920 | n4005 ;
  assign n11525 = x[73] & n3906 ;
  assign n11526 = n11524 | n11525 ;
  assign n11527 = n4044 | n11526 ;
  assign n29332 = ~n11527 ;
  assign n11528 = x[35] & n29332 ;
  assign n11529 = n28822 & n11527 ;
  assign n11530 = n11528 | n11529 ;
  assign n11531 = n11523 & n11530 ;
  assign n11643 = n11523 | n11530 ;
  assign n29333 = ~n11531 ;
  assign n12145 = n29333 & n11643 ;
  assign n12146 = n11642 & n12145 ;
  assign n12464 = n11642 | n12145 ;
  assign n29334 = ~n12146 ;
  assign n12465 = n29334 & n12464 ;
  assign n29335 = ~n12311 ;
  assign n12467 = n29335 & n12465 ;
  assign n29336 = ~n12465 ;
  assign n12865 = n12311 & n29336 ;
  assign n12866 = n12467 | n12865 ;
  assign n12867 = n12463 | n12866 ;
  assign n12869 = n12463 & n12866 ;
  assign n29337 = ~n12869 ;
  assign n13177 = n12867 & n29337 ;
  assign n4635 = n1741 & n4632 ;
  assign n4548 = x[77] & n4514 ;
  assign n4620 = x[78] & n4572 ;
  assign n13178 = n4548 | n4620 ;
  assign n13179 = x[79] & n4504 ;
  assign n13180 = n13178 | n13179 ;
  assign n13181 = n4635 | n13180 ;
  assign n29338 = ~n13181 ;
  assign n13182 = x[29] & n29338 ;
  assign n13183 = n28483 & n13181 ;
  assign n13184 = n13182 | n13183 ;
  assign n29339 = ~n13184 ;
  assign n13185 = n13177 & n29339 ;
  assign n29340 = ~n13177 ;
  assign n13785 = n29340 & n13184 ;
  assign n13786 = n13185 | n13785 ;
  assign n29341 = ~n13786 ;
  assign n13787 = n13385 & n29341 ;
  assign n29342 = ~n13385 ;
  assign n13915 = n29342 & n13786 ;
  assign n13916 = n13787 | n13915 ;
  assign n1004 = n452 & n1003 ;
  assign n386 = x[80] & n330 ;
  assign n397 = x[81] & n390 ;
  assign n13917 = n386 | n397 ;
  assign n13918 = x[82] & n322 ;
  assign n13919 = n13917 | n13918 ;
  assign n13920 = n1004 | n13919 ;
  assign n29343 = ~n13920 ;
  assign n13921 = x[26] & n29343 ;
  assign n13922 = n28342 & n13920 ;
  assign n13923 = n13921 | n13922 ;
  assign n13924 = n13916 | n13923 ;
  assign n13925 = n13916 & n13923 ;
  assign n29344 = ~n13925 ;
  assign n14734 = n13924 & n29344 ;
  assign n29345 = ~n14176 ;
  assign n14736 = n29345 & n14734 ;
  assign n29346 = ~n14734 ;
  assign n14821 = n14176 & n29346 ;
  assign n14822 = n14736 | n14821 ;
  assign n14823 = n14820 & n14822 ;
  assign n14825 = n14820 | n14822 ;
  assign n29347 = ~n14823 ;
  assign n14826 = n29347 & n14825 ;
  assign n15790 = n14853 | n15789 ;
  assign n15791 = n15730 & n15790 ;
  assign n15792 = n14836 | n15791 ;
  assign n29348 = ~n15792 ;
  assign n15793 = n14826 & n29348 ;
  assign n29349 = ~n14826 ;
  assign n15829 = n29349 & n15792 ;
  assign n15830 = n15793 | n15829 ;
  assign n7176 = n1720 & n7162 ;
  assign n7113 = x[86] & n7100 ;
  assign n7699 = x[87] & n7647 ;
  assign n15831 = n7113 | n7699 ;
  assign n15832 = x[88] & n7098 ;
  assign n15833 = n15831 | n15832 ;
  assign n15834 = n7176 | n15833 ;
  assign n29350 = ~n15834 ;
  assign n15835 = x[20] & n29350 ;
  assign n15836 = n28114 & n15834 ;
  assign n15837 = n15835 | n15836 ;
  assign n15838 = n15830 & n15837 ;
  assign n29351 = ~n14820 ;
  assign n14824 = n29351 & n14822 ;
  assign n29352 = ~n14822 ;
  assign n15727 = n14820 & n29352 ;
  assign n15728 = n14824 | n15727 ;
  assign n15794 = n15728 | n15792 ;
  assign n15795 = n15728 & n15792 ;
  assign n29353 = ~n15795 ;
  assign n16173 = n15794 & n29353 ;
  assign n16174 = n15837 | n16173 ;
  assign n29354 = ~n15838 ;
  assign n16476 = n29354 & n16174 ;
  assign n29355 = ~n16172 ;
  assign n16478 = n29355 & n16476 ;
  assign n29356 = ~n16476 ;
  assign n16747 = n16172 & n29356 ;
  assign n16748 = n16478 | n16747 ;
  assign n29357 = ~n16746 ;
  assign n17133 = n29357 & n16748 ;
  assign n29358 = ~n16748 ;
  assign n17464 = n16746 & n29358 ;
  assign n17465 = n17133 | n17464 ;
  assign n17466 = n17463 | n17465 ;
  assign n17467 = n17463 & n17465 ;
  assign n29359 = ~n17467 ;
  assign n17708 = n17466 & n29359 ;
  assign n10568 = n2410 & n10542 ;
  assign n10508 = x[92] & n10481 ;
  assign n11884 = x[93] & n11232 ;
  assign n17709 = n10508 | n11884 ;
  assign n17710 = x[94] & n10479 ;
  assign n17711 = n17709 | n17710 ;
  assign n17712 = n10568 | n17711 ;
  assign n29360 = ~n17712 ;
  assign n17713 = x[14] & n29360 ;
  assign n17714 = n27956 & n17712 ;
  assign n17715 = n17713 | n17714 ;
  assign n17716 = n17708 | n17715 ;
  assign n17717 = n17708 & n17715 ;
  assign n29361 = ~n17717 ;
  assign n18732 = n17716 & n29361 ;
  assign n29362 = ~n18216 ;
  assign n18734 = n29362 & n18732 ;
  assign n29363 = ~n18732 ;
  assign n18964 = n18216 & n29363 ;
  assign n18965 = n18734 | n18964 ;
  assign n29364 = ~n18963 ;
  assign n19510 = n29364 & n18965 ;
  assign n29365 = ~n18965 ;
  assign n19511 = n18963 & n29365 ;
  assign n19512 = n19510 | n19511 ;
  assign n19513 = n19509 | n19512 ;
  assign n19514 = n19509 & n19512 ;
  assign n29366 = ~n19514 ;
  assign n20235 = n19513 & n29366 ;
  assign n15357 = n2466 & n15308 ;
  assign n15305 = x[98] & n15246 ;
  assign n17318 = x[99] & n16288 ;
  assign n20236 = n15305 | n17318 ;
  assign n20237 = x[100] & n15244 ;
  assign n20238 = n20236 | n20237 ;
  assign n20239 = n15357 | n20238 ;
  assign n29367 = ~n20239 ;
  assign n20240 = x[8] & n29367 ;
  assign n20241 = n27845 & n20239 ;
  assign n20242 = n20240 | n20241 ;
  assign n20243 = n20235 | n20242 ;
  assign n20244 = n20235 & n20242 ;
  assign n29368 = ~n20244 ;
  assign n21266 = n20243 & n29368 ;
  assign n21267 = n21265 & n21266 ;
  assign n21977 = n21265 | n21266 ;
  assign n29369 = ~n21267 ;
  assign n21978 = n29369 & n21977 ;
  assign n29370 = ~n21403 ;
  assign n21980 = n29370 & n21978 ;
  assign n29371 = ~n21978 ;
  assign n22265 = n21403 & n29371 ;
  assign n22266 = n21980 | n22265 ;
  assign n22267 = n22264 | n22266 ;
  assign n22268 = n22264 & n22266 ;
  assign n29372 = ~n22268 ;
  assign n22403 = n22267 & n29372 ;
  assign n579 = n577 & n578 ;
  assign n580 = n27622 | n579 ;
  assign n25068 = x[105] & x[106] ;
  assign n581 = x[105] | x[106] ;
  assign n29373 = ~n25068 ;
  assign n3220 = n29373 & n581 ;
  assign n3221 = n580 & n3220 ;
  assign n3222 = n580 | n3220 ;
  assign n29374 = ~n3221 ;
  assign n3223 = n29374 & n3222 ;
  assign n19714 = n3223 & n19656 ;
  assign n19777 = x[104] & n19723 ;
  assign n19880 = x[105] & n19829 ;
  assign n22404 = n19777 | n19880 ;
  assign n22405 = x[106] & n19655 ;
  assign n22406 = n22404 | n22405 ;
  assign n22407 = n19714 | n22406 ;
  assign n29375 = ~n22407 ;
  assign n22408 = x[2] & n29375 ;
  assign n22409 = n27790 & n22407 ;
  assign n22410 = n22408 | n22409 ;
  assign n29376 = ~n22410 ;
  assign n22411 = n22403 & n29376 ;
  assign n29377 = ~n22403 ;
  assign n22413 = n29377 & n22410 ;
  assign n22414 = n22411 | n22413 ;
  assign n23013 = n22425 | n23012 ;
  assign n23014 = n22414 & n23013 ;
  assign n27684 = n22414 | n23013 ;
  assign n29378 = ~n23014 ;
  assign n171 = n29378 & n27684 ;
  assign n582 = n580 & n581 ;
  assign n583 = n25068 | n582 ;
  assign n27620 = x[106] & x[107] ;
  assign n584 = x[106] | x[107] ;
  assign n29379 = ~n27620 ;
  assign n3196 = n29379 & n584 ;
  assign n29380 = ~n583 ;
  assign n3197 = n29380 & n3196 ;
  assign n29381 = ~n3196 ;
  assign n3198 = n583 & n29381 ;
  assign n3199 = n3197 | n3198 ;
  assign n19711 = n3199 & n19656 ;
  assign n19762 = x[105] & n19723 ;
  assign n19881 = x[106] & n19829 ;
  assign n22391 = n19762 | n19881 ;
  assign n22392 = x[107] & n19655 ;
  assign n22393 = n22391 | n22392 ;
  assign n22394 = n19711 | n22393 ;
  assign n29382 = ~n22394 ;
  assign n22395 = x[2] & n29382 ;
  assign n22396 = n27790 & n22394 ;
  assign n22397 = n22395 | n22396 ;
  assign n20851 = n20251 | n20253 ;
  assign n29383 = ~n20254 ;
  assign n20852 = n29383 & n20851 ;
  assign n20853 = n20849 & n20852 ;
  assign n20854 = n20254 | n20853 ;
  assign n29384 = ~n20854 ;
  assign n21268 = n29384 & n21266 ;
  assign n29385 = ~n21266 ;
  assign n21404 = n20854 & n29385 ;
  assign n21405 = n21268 | n21404 ;
  assign n21406 = n21403 & n21405 ;
  assign n22269 = n21406 | n22268 ;
  assign n12720 = n2841 & n12695 ;
  assign n12664 = x[96] & n12633 ;
  assign n14408 = x[97] & n13533 ;
  assign n18944 = n12664 | n14408 ;
  assign n18945 = x[98] & n12631 ;
  assign n18946 = n18944 | n18945 ;
  assign n18947 = n12720 | n18946 ;
  assign n29386 = ~n18947 ;
  assign n18948 = x[11] & n29386 ;
  assign n18949 = n27892 & n18947 ;
  assign n18950 = n18948 | n18949 ;
  assign n8727 = n1841 & n8706 ;
  assign n8652 = x[90] & n8645 ;
  assign n9885 = x[91] & n9278 ;
  assign n16730 = n8652 | n9885 ;
  assign n16731 = x[92] & n8643 ;
  assign n16732 = n16730 | n16731 ;
  assign n16733 = n8727 | n16732 ;
  assign n29387 = ~n16733 ;
  assign n16734 = x[17] & n29387 ;
  assign n16735 = n28039 & n16733 ;
  assign n16736 = n16734 | n16735 ;
  assign n5313 = n1213 & n5302 ;
  assign n5251 = x[84] & n5240 ;
  assign n6234 = x[85] & n6179 ;
  assign n14801 = n5251 | n6234 ;
  assign n14802 = x[86] & n5238 ;
  assign n14803 = n14801 | n14802 ;
  assign n14804 = n5313 | n14803 ;
  assign n29388 = ~n14804 ;
  assign n14805 = x[23] & n29388 ;
  assign n14806 = n28221 & n14804 ;
  assign n14807 = n14805 | n14806 ;
  assign n4642 = n1270 & n4632 ;
  assign n4561 = x[78] & n4514 ;
  assign n4619 = x[79] & n4572 ;
  assign n13164 = n4561 | n4619 ;
  assign n13165 = x[80] & n4504 ;
  assign n13166 = n13164 | n13165 ;
  assign n13167 = n4642 | n13166 ;
  assign n29389 = ~n13167 ;
  assign n13168 = x[29] & n29389 ;
  assign n13169 = n28483 & n13167 ;
  assign n13170 = n13168 | n13169 ;
  assign n29390 = ~n11642 ;
  assign n12147 = n29390 & n12145 ;
  assign n29391 = ~n12145 ;
  assign n12312 = n11642 & n29391 ;
  assign n12313 = n12147 | n12312 ;
  assign n12314 = n12311 & n12313 ;
  assign n12870 = n12314 | n12869 ;
  assign n4798 = n3574 & n4790 ;
  assign n3486 = x[69] & n3443 ;
  assign n3524 = x[70] & n3508 ;
  assign n10946 = n3486 | n3524 ;
  assign n10947 = x[71] & n3439 ;
  assign n10948 = n10946 | n10947 ;
  assign n10949 = n4798 | n10948 ;
  assign n29392 = ~n10949 ;
  assign n10950 = x[38] & n29392 ;
  assign n10951 = n28996 & n10949 ;
  assign n10952 = n10950 | n10951 ;
  assign n10270 = n10261 & n10268 ;
  assign n10271 = n10259 | n10270 ;
  assign n6411 = n3162 & n6408 ;
  assign n3042 = x[66] & n3031 ;
  assign n3113 = x[67] & n3096 ;
  assign n10229 = n3042 | n3113 ;
  assign n10230 = x[68] & n3027 ;
  assign n10231 = n10229 | n10230 ;
  assign n10232 = n6411 | n10231 ;
  assign n10233 = x[41] | n10232 ;
  assign n10234 = x[41] & n10232 ;
  assign n29393 = ~n10234 ;
  assign n10235 = n10233 & n29393 ;
  assign n29394 = ~n9557 ;
  assign n9558 = x[44] & n29394 ;
  assign n27707 = x[43] & x[44] ;
  assign n2486 = x[43] | x[44] ;
  assign n29395 = ~n27707 ;
  assign n2487 = n29395 & n2486 ;
  assign n2635 = n2485 & n2487 ;
  assign n6440 = n2635 & n6437 ;
  assign n29396 = ~n2487 ;
  assign n2488 = n2485 & n29396 ;
  assign n9559 = x[65] & n2488 ;
  assign n27709 = x[42] & x[43] ;
  assign n2489 = x[42] | x[43] ;
  assign n29397 = ~n27709 ;
  assign n2490 = n29397 & n2489 ;
  assign n29398 = ~n2485 ;
  assign n2557 = n29398 & n2490 ;
  assign n9560 = x[64] & n2557 ;
  assign n9561 = n9559 | n9560 ;
  assign n9562 = n6440 | n9561 ;
  assign n29399 = ~n9562 ;
  assign n9563 = x[44] & n29399 ;
  assign n29400 = ~x[44] ;
  assign n9564 = n29400 & n9562 ;
  assign n9565 = n9563 | n9564 ;
  assign n29401 = ~n9565 ;
  assign n9566 = n9558 & n29401 ;
  assign n29402 = ~n9558 ;
  assign n10236 = n29402 & n9565 ;
  assign n10237 = n9566 | n10236 ;
  assign n10238 = n10235 & n10237 ;
  assign n10272 = n10235 | n10237 ;
  assign n29403 = ~n10238 ;
  assign n10273 = n29403 & n10272 ;
  assign n29404 = ~n10271 ;
  assign n10274 = n29404 & n10273 ;
  assign n29405 = ~n10273 ;
  assign n10953 = n10271 & n29405 ;
  assign n10954 = n10274 | n10953 ;
  assign n29406 = ~n10952 ;
  assign n10955 = n29406 & n10954 ;
  assign n29407 = ~n10954 ;
  assign n10957 = n10952 & n29407 ;
  assign n10958 = n10955 | n10957 ;
  assign n11036 = n10970 & n11034 ;
  assign n11037 = n10968 | n11036 ;
  assign n29408 = ~n11037 ;
  assign n11038 = n10958 & n29408 ;
  assign n29409 = ~n10958 ;
  assign n11512 = n29409 & n11037 ;
  assign n11513 = n11038 | n11512 ;
  assign n4045 = n2722 & n4041 ;
  assign n3954 = x[72] & n3910 ;
  assign n3984 = x[73] & n3975 ;
  assign n11514 = n3954 | n3984 ;
  assign n11515 = x[74] & n3906 ;
  assign n11516 = n11514 | n11515 ;
  assign n11517 = n4045 | n11516 ;
  assign n29410 = ~n11517 ;
  assign n11518 = x[35] & n29410 ;
  assign n11519 = n28822 & n11517 ;
  assign n11520 = n11518 | n11519 ;
  assign n11646 = n11513 | n11520 ;
  assign n11521 = n11513 & n11520 ;
  assign n11644 = n11642 & n11643 ;
  assign n11645 = n11531 | n11644 ;
  assign n11647 = n11645 & n11646 ;
  assign n11649 = n11521 | n11647 ;
  assign n29411 = ~n11649 ;
  assign n11650 = n11646 & n29411 ;
  assign n29412 = ~n11521 ;
  assign n11648 = n29412 & n11646 ;
  assign n12148 = n11531 | n12146 ;
  assign n29413 = ~n11648 ;
  assign n12294 = n29413 & n12148 ;
  assign n12295 = n11650 | n12294 ;
  assign n1777 = n779 & n1775 ;
  assign n713 = x[75] & n663 ;
  assign n765 = x[76] & n720 ;
  assign n12296 = n713 | n765 ;
  assign n12297 = x[77] & n652 ;
  assign n12298 = n12296 | n12297 ;
  assign n12299 = n1777 | n12298 ;
  assign n29414 = ~n12299 ;
  assign n12300 = x[32] & n29414 ;
  assign n12301 = n28658 & n12299 ;
  assign n12302 = n12300 | n12301 ;
  assign n12303 = n12295 | n12302 ;
  assign n12304 = n12295 & n12302 ;
  assign n29415 = ~n12304 ;
  assign n12871 = n12303 & n29415 ;
  assign n12872 = n12870 & n12871 ;
  assign n13171 = n12870 | n12871 ;
  assign n29416 = ~n12872 ;
  assign n13172 = n29416 & n13171 ;
  assign n29417 = ~n13170 ;
  assign n13174 = n29417 & n13172 ;
  assign n29418 = ~n13172 ;
  assign n13175 = n13170 & n29418 ;
  assign n13176 = n13174 | n13175 ;
  assign n13186 = n13177 & n13184 ;
  assign n29419 = ~n12866 ;
  assign n12868 = n12463 & n29419 ;
  assign n29420 = ~n12463 ;
  assign n13386 = n29420 & n12866 ;
  assign n13387 = n12868 | n13386 ;
  assign n13388 = n13184 | n13387 ;
  assign n13389 = n13184 & n13387 ;
  assign n29421 = ~n13389 ;
  assign n13390 = n13388 & n29421 ;
  assign n13391 = n13385 & n13390 ;
  assign n13392 = n13186 | n13391 ;
  assign n13393 = n13176 | n13392 ;
  assign n13394 = n13176 & n13392 ;
  assign n29422 = ~n13394 ;
  assign n13900 = n13393 & n29422 ;
  assign n1059 = n452 & n1057 ;
  assign n343 = x[81] & n330 ;
  assign n440 = x[82] & n390 ;
  assign n13901 = n343 | n440 ;
  assign n13902 = x[83] & n322 ;
  assign n13903 = n13901 | n13902 ;
  assign n13904 = n1059 | n13903 ;
  assign n29423 = ~n13904 ;
  assign n13905 = x[26] & n29423 ;
  assign n13906 = n28342 & n13904 ;
  assign n13907 = n13905 | n13906 ;
  assign n29424 = ~n13907 ;
  assign n13908 = n13900 & n29424 ;
  assign n29425 = ~n13900 ;
  assign n14696 = n29425 & n13907 ;
  assign n14697 = n13908 | n14696 ;
  assign n14729 = n13958 | n14728 ;
  assign n14730 = n14699 & n14729 ;
  assign n14731 = n13945 | n14730 ;
  assign n14732 = n14173 & n14731 ;
  assign n14733 = n13935 | n14732 ;
  assign n14735 = n14733 & n14734 ;
  assign n14737 = n13925 | n14735 ;
  assign n14739 = n14697 | n14737 ;
  assign n14740 = n14697 & n14737 ;
  assign n29426 = ~n14740 ;
  assign n14810 = n14739 & n29426 ;
  assign n29427 = ~n14807 ;
  assign n14811 = n29427 & n14810 ;
  assign n29428 = ~n14810 ;
  assign n14812 = n14807 & n29428 ;
  assign n14813 = n14811 | n14812 ;
  assign n15111 = n14836 | n15110 ;
  assign n15112 = n14826 & n15111 ;
  assign n15113 = n14823 | n15112 ;
  assign n15114 = n14813 | n15113 ;
  assign n15115 = n14813 & n15113 ;
  assign n29429 = ~n15115 ;
  assign n15814 = n15114 & n29429 ;
  assign n7170 = n1453 & n7162 ;
  assign n7138 = x[87] & n7100 ;
  assign n7687 = x[88] & n7647 ;
  assign n15815 = n7138 | n7687 ;
  assign n15816 = x[89] & n7098 ;
  assign n15817 = n15815 | n15816 ;
  assign n15818 = n7170 | n15817 ;
  assign n29430 = ~n15818 ;
  assign n15819 = x[20] & n29430 ;
  assign n15820 = n28114 & n15818 ;
  assign n15821 = n15819 | n15820 ;
  assign n29431 = ~n15821 ;
  assign n15822 = n15814 & n29431 ;
  assign n29432 = ~n15814 ;
  assign n16402 = n29432 & n15821 ;
  assign n16403 = n15822 | n16402 ;
  assign n16404 = n15837 & n16173 ;
  assign n16477 = n16475 & n16476 ;
  assign n16479 = n16404 | n16477 ;
  assign n16481 = n16403 | n16479 ;
  assign n16482 = n16403 & n16479 ;
  assign n29433 = ~n16482 ;
  assign n17138 = n16481 & n29433 ;
  assign n29434 = ~n16736 ;
  assign n17139 = n29434 & n17138 ;
  assign n29435 = ~n17138 ;
  assign n17141 = n16736 & n29435 ;
  assign n17142 = n17139 | n17141 ;
  assign n16749 = n16746 & n16748 ;
  assign n17468 = n16749 | n17467 ;
  assign n29436 = ~n17142 ;
  assign n17469 = n29436 & n17468 ;
  assign n29437 = ~n17468 ;
  assign n17698 = n17142 & n29437 ;
  assign n17699 = n17469 | n17698 ;
  assign n10602 = n2152 & n10542 ;
  assign n10507 = x[93] & n10481 ;
  assign n11908 = x[94] & n11232 ;
  assign n17700 = n10507 | n11908 ;
  assign n17701 = x[95] & n10479 ;
  assign n17702 = n17700 | n17701 ;
  assign n17703 = n10602 | n17702 ;
  assign n29438 = ~n17703 ;
  assign n17704 = x[14] & n29438 ;
  assign n17705 = n27956 & n17703 ;
  assign n17706 = n17704 | n17705 ;
  assign n17707 = n17699 & n17706 ;
  assign n18219 = n17699 | n17706 ;
  assign n29439 = ~n17707 ;
  assign n18220 = n29439 & n18219 ;
  assign n18208 = n17734 & n18206 ;
  assign n18726 = n17734 | n18206 ;
  assign n29440 = ~n18208 ;
  assign n18727 = n29440 & n18726 ;
  assign n18728 = n18724 & n18727 ;
  assign n18729 = n17737 | n18728 ;
  assign n18730 = n18213 & n18729 ;
  assign n18731 = n17727 | n18730 ;
  assign n18733 = n18731 & n18732 ;
  assign n18735 = n17717 | n18733 ;
  assign n29441 = ~n18735 ;
  assign n18736 = n18220 & n29441 ;
  assign n29442 = ~n18220 ;
  assign n18951 = n29442 & n18735 ;
  assign n18952 = n18736 | n18951 ;
  assign n29443 = ~n18950 ;
  assign n18954 = n29443 & n18952 ;
  assign n29444 = ~n18952 ;
  assign n20058 = n18950 & n29444 ;
  assign n20059 = n18954 | n20058 ;
  assign n18966 = n18963 & n18965 ;
  assign n20080 = n19506 & n20078 ;
  assign n20081 = n18976 | n20080 ;
  assign n20082 = n18963 | n18965 ;
  assign n29445 = ~n18966 ;
  assign n20083 = n29445 & n20082 ;
  assign n20084 = n20081 & n20083 ;
  assign n20085 = n18966 | n20084 ;
  assign n20086 = n20059 | n20085 ;
  assign n20088 = n20059 & n20085 ;
  assign n29446 = ~n20088 ;
  assign n20226 = n20086 & n29446 ;
  assign n15355 = n2977 & n15308 ;
  assign n15272 = x[99] & n15246 ;
  assign n17322 = x[100] & n16288 ;
  assign n20227 = n15272 | n17322 ;
  assign n20228 = x[101] & n15244 ;
  assign n20229 = n20227 | n20228 ;
  assign n20230 = n15355 | n20229 ;
  assign n29447 = ~n20230 ;
  assign n20231 = x[8] & n29447 ;
  assign n20232 = n27845 & n20230 ;
  assign n20233 = n20231 | n20232 ;
  assign n20857 = n20226 | n20233 ;
  assign n20234 = n20226 & n20233 ;
  assign n20855 = n20243 & n20854 ;
  assign n20856 = n20244 | n20855 ;
  assign n20858 = n20856 & n20857 ;
  assign n20859 = n20234 | n20858 ;
  assign n29448 = ~n20859 ;
  assign n20860 = n20857 & n29448 ;
  assign n18953 = n18950 & n18952 ;
  assign n18955 = n18950 | n18952 ;
  assign n29449 = ~n18953 ;
  assign n18956 = n29449 & n18955 ;
  assign n29450 = ~n20085 ;
  assign n20087 = n18956 & n29450 ;
  assign n29451 = ~n18956 ;
  assign n21118 = n29451 & n20085 ;
  assign n21119 = n20087 | n21118 ;
  assign n21120 = n20233 & n21119 ;
  assign n29452 = ~n21120 ;
  assign n21121 = n20857 & n29452 ;
  assign n21269 = n20244 | n21267 ;
  assign n29453 = ~n21121 ;
  assign n21386 = n29453 & n21269 ;
  assign n21387 = n20860 | n21386 ;
  assign n18452 = n3001 & n18392 ;
  assign n18383 = x[102] & n18329 ;
  assign n18526 = x[103] & n18514 ;
  assign n21388 = n18383 | n18526 ;
  assign n21389 = x[104] & n18327 ;
  assign n21390 = n21388 | n21389 ;
  assign n21391 = n18452 | n21390 ;
  assign n29454 = ~n21391 ;
  assign n21392 = x[5] & n29454 ;
  assign n21393 = n27813 & n21391 ;
  assign n21394 = n21392 | n21393 ;
  assign n21395 = n21387 | n21394 ;
  assign n21396 = n21387 & n21394 ;
  assign n29455 = ~n21396 ;
  assign n22270 = n21395 & n29455 ;
  assign n22271 = n22269 & n22270 ;
  assign n22398 = n22269 | n22270 ;
  assign n29456 = ~n22271 ;
  assign n22399 = n29456 & n22398 ;
  assign n22400 = n22397 | n22399 ;
  assign n22401 = n22397 & n22399 ;
  assign n29457 = ~n22401 ;
  assign n22402 = n22400 & n29457 ;
  assign n22412 = n22403 & n22410 ;
  assign n23015 = n22412 | n23014 ;
  assign n23016 = n22402 | n23015 ;
  assign n23017 = n22402 & n23015 ;
  assign n29458 = ~n23017 ;
  assign n172 = n23016 & n29458 ;
  assign n23018 = n22401 | n23017 ;
  assign n22272 = n21396 | n22271 ;
  assign n18434 = n3409 & n18392 ;
  assign n18365 = x[103] & n18329 ;
  assign n18572 = x[104] & n18514 ;
  assign n21376 = n18365 | n18572 ;
  assign n21377 = x[105] & n18327 ;
  assign n21378 = n21376 | n21377 ;
  assign n21379 = n18434 | n21378 ;
  assign n29459 = ~n21379 ;
  assign n21380 = x[5] & n29459 ;
  assign n21381 = n27813 & n21379 ;
  assign n21382 = n21380 | n21381 ;
  assign n15361 = n2867 & n15308 ;
  assign n15302 = x[100] & n15246 ;
  assign n17308 = x[101] & n16288 ;
  assign n20217 = n15302 | n17308 ;
  assign n20218 = x[102] & n15244 ;
  assign n20219 = n20217 | n20218 ;
  assign n20220 = n15361 | n20219 ;
  assign n29460 = ~n20220 ;
  assign n20221 = x[8] & n29460 ;
  assign n20222 = n27845 & n20220 ;
  assign n20223 = n20221 | n20222 ;
  assign n12721 = n2313 & n12695 ;
  assign n12666 = x[97] & n12633 ;
  assign n14407 = x[98] & n13533 ;
  assign n18931 = n12666 | n14407 ;
  assign n18932 = x[99] & n12631 ;
  assign n18933 = n18931 | n18932 ;
  assign n18934 = n12721 | n18933 ;
  assign n29461 = ~n18934 ;
  assign n18935 = x[11] & n29461 ;
  assign n18936 = n27892 & n18934 ;
  assign n18937 = n18935 | n18936 ;
  assign n18217 = n17716 & n18216 ;
  assign n18218 = n17717 | n18217 ;
  assign n18221 = n18218 & n18220 ;
  assign n18222 = n17707 | n18221 ;
  assign n10566 = n2000 & n10542 ;
  assign n10510 = x[94] & n10481 ;
  assign n11876 = x[95] & n11232 ;
  assign n17688 = n10510 | n11876 ;
  assign n17689 = x[96] & n10479 ;
  assign n17690 = n17688 | n17689 ;
  assign n17691 = n10566 | n17690 ;
  assign n29462 = ~n17691 ;
  assign n17692 = x[14] & n29462 ;
  assign n17693 = n27956 & n17691 ;
  assign n17694 = n17692 | n17693 ;
  assign n13173 = n13170 & n13172 ;
  assign n13763 = n13170 | n13172 ;
  assign n29463 = ~n13173 ;
  assign n13764 = n29463 & n13763 ;
  assign n29464 = ~n13392 ;
  assign n13765 = n29464 & n13764 ;
  assign n29465 = ~n13764 ;
  assign n13910 = n13392 & n29465 ;
  assign n13911 = n13765 | n13910 ;
  assign n13912 = n13907 | n13911 ;
  assign n13913 = n13907 & n13911 ;
  assign n29466 = ~n13913 ;
  assign n13914 = n13912 & n29466 ;
  assign n29467 = ~n14737 ;
  assign n14738 = n13914 & n29467 ;
  assign n29468 = ~n13914 ;
  assign n14799 = n29468 & n14737 ;
  assign n14800 = n14738 | n14799 ;
  assign n14808 = n14800 | n14807 ;
  assign n14809 = n14800 & n14807 ;
  assign n29469 = ~n14809 ;
  assign n15725 = n14808 & n29469 ;
  assign n29470 = ~n15113 ;
  assign n15726 = n29470 & n15725 ;
  assign n29471 = ~n15725 ;
  assign n15824 = n15113 & n29471 ;
  assign n15825 = n15726 | n15824 ;
  assign n15826 = n15821 | n15825 ;
  assign n15827 = n15821 & n15825 ;
  assign n29472 = ~n15827 ;
  assign n15828 = n15826 & n29472 ;
  assign n29473 = ~n16479 ;
  assign n16480 = n15828 & n29473 ;
  assign n29474 = ~n15828 ;
  assign n16737 = n29474 & n16479 ;
  assign n16738 = n16480 | n16737 ;
  assign n16739 = n16736 & n16738 ;
  assign n16772 = n16763 & n16770 ;
  assign n17128 = n16777 & n17127 ;
  assign n17129 = n16772 | n17128 ;
  assign n17130 = n16753 | n16760 ;
  assign n17131 = n17129 & n17130 ;
  assign n17132 = n16762 | n17131 ;
  assign n17134 = n16746 | n16748 ;
  assign n29475 = ~n16749 ;
  assign n17135 = n29475 & n17134 ;
  assign n17136 = n17132 & n17135 ;
  assign n17137 = n16749 | n17136 ;
  assign n17143 = n17137 & n17142 ;
  assign n17144 = n16739 | n17143 ;
  assign n8735 = n1685 & n8706 ;
  assign n8673 = x[91] & n8645 ;
  assign n9883 = x[92] & n9278 ;
  assign n16720 = n8673 | n9883 ;
  assign n16721 = x[93] & n8643 ;
  assign n16722 = n16720 | n16721 ;
  assign n16723 = n8735 | n16722 ;
  assign n29476 = ~n16723 ;
  assign n16724 = x[17] & n29476 ;
  assign n16725 = n28039 & n16723 ;
  assign n16726 = n16724 | n16725 ;
  assign n16483 = n15827 | n16482 ;
  assign n15116 = n14809 | n15115 ;
  assign n1294 = n452 & n1293 ;
  assign n344 = x[82] & n330 ;
  assign n439 = x[83] & n390 ;
  assign n13887 = n344 | n439 ;
  assign n13888 = x[84] & n322 ;
  assign n13889 = n13887 | n13888 ;
  assign n13890 = n1294 | n13889 ;
  assign n29477 = ~n13890 ;
  assign n13891 = x[26] & n29477 ;
  assign n13892 = n28342 & n13890 ;
  assign n13893 = n13891 | n13892 ;
  assign n13395 = n13173 | n13394 ;
  assign n4638 = n1029 & n4632 ;
  assign n4556 = x[79] & n4514 ;
  assign n4598 = x[80] & n4572 ;
  assign n13154 = n4556 | n4598 ;
  assign n13155 = x[81] & n4504 ;
  assign n13156 = n13154 | n13155 ;
  assign n13157 = n4638 | n13156 ;
  assign n29478 = ~n13157 ;
  assign n13158 = x[29] & n29478 ;
  assign n13159 = n28483 & n13157 ;
  assign n13160 = n13158 | n13159 ;
  assign n2086 = n779 & n2084 ;
  assign n712 = x[76] & n663 ;
  assign n764 = x[77] & n720 ;
  assign n12284 = n712 | n764 ;
  assign n12285 = x[78] & n652 ;
  assign n12286 = n12284 | n12285 ;
  assign n12287 = n2086 | n12286 ;
  assign n29479 = ~n12287 ;
  assign n12288 = x[32] & n29479 ;
  assign n12289 = n28658 & n12287 ;
  assign n12290 = n12288 | n12289 ;
  assign n12149 = n11646 & n12148 ;
  assign n12150 = n11521 | n12149 ;
  assign n10956 = n10952 & n10954 ;
  assign n11039 = n10958 & n11037 ;
  assign n11040 = n10956 | n11039 ;
  assign n3704 = n3574 & n3701 ;
  assign n3463 = x[70] & n3443 ;
  assign n3517 = x[71] & n3508 ;
  assign n10935 = n3463 | n3517 ;
  assign n10936 = x[72] & n3439 ;
  assign n10937 = n10935 | n10936 ;
  assign n10938 = n3704 | n10937 ;
  assign n29480 = ~n10938 ;
  assign n10939 = x[38] & n29480 ;
  assign n10940 = n28996 & n10938 ;
  assign n10941 = n10939 | n10940 ;
  assign n10275 = n10271 & n10273 ;
  assign n10276 = n10238 | n10275 ;
  assign n9567 = n9558 & n9565 ;
  assign n6471 = n2635 & n6466 ;
  assign n2491 = n29398 & n2487 ;
  assign n29481 = ~n2490 ;
  assign n2492 = n29481 & n2491 ;
  assign n2500 = x[64] & n2492 ;
  assign n2569 = x[65] & n2557 ;
  assign n9568 = n2500 | n2569 ;
  assign n9569 = x[66] & n2488 ;
  assign n9570 = n9568 | n9569 ;
  assign n9571 = n6471 | n9570 ;
  assign n29482 = ~n9571 ;
  assign n9572 = x[44] & n29482 ;
  assign n9573 = n29400 & n9571 ;
  assign n9574 = n9572 | n9573 ;
  assign n29483 = ~n9574 ;
  assign n9575 = n9567 & n29483 ;
  assign n29484 = ~n9567 ;
  assign n10218 = n29484 & n9574 ;
  assign n10219 = n9575 | n10218 ;
  assign n6388 = n3162 & n6379 ;
  assign n3063 = x[67] & n3031 ;
  assign n3114 = x[68] & n3096 ;
  assign n10220 = n3063 | n3114 ;
  assign n10221 = x[69] & n3027 ;
  assign n10222 = n10220 | n10221 ;
  assign n10223 = n6388 | n10222 ;
  assign n29485 = ~n10223 ;
  assign n10224 = x[41] & n29485 ;
  assign n10225 = n29184 & n10223 ;
  assign n10226 = n10224 | n10225 ;
  assign n29486 = ~n10226 ;
  assign n10227 = n10219 & n29486 ;
  assign n29487 = ~n10219 ;
  assign n10277 = n29487 & n10226 ;
  assign n10278 = n10227 | n10277 ;
  assign n29488 = ~n10278 ;
  assign n10279 = n10276 & n29488 ;
  assign n29489 = ~n10276 ;
  assign n10942 = n29489 & n10278 ;
  assign n10943 = n10279 | n10942 ;
  assign n29490 = ~n10941 ;
  assign n10944 = n29490 & n10943 ;
  assign n29491 = ~n10943 ;
  assign n11041 = n10941 & n29491 ;
  assign n11042 = n10944 | n11041 ;
  assign n29492 = ~n11042 ;
  assign n11475 = n11040 & n29492 ;
  assign n29493 = ~n11040 ;
  assign n11502 = n29493 & n11042 ;
  assign n11503 = n11475 | n11502 ;
  assign n4068 = n3289 & n4041 ;
  assign n3925 = x[73] & n3910 ;
  assign n3986 = x[74] & n3975 ;
  assign n11504 = n3925 | n3986 ;
  assign n11505 = x[75] & n3906 ;
  assign n11506 = n11504 | n11505 ;
  assign n11507 = n4068 | n11506 ;
  assign n29494 = ~n11507 ;
  assign n11508 = x[35] & n29494 ;
  assign n11509 = n28822 & n11507 ;
  assign n11510 = n11508 | n11509 ;
  assign n11511 = n11503 & n11510 ;
  assign n11043 = n11040 | n11042 ;
  assign n11044 = n11040 & n11042 ;
  assign n29495 = ~n11044 ;
  assign n11651 = n11043 & n29495 ;
  assign n11652 = n11510 | n11651 ;
  assign n29496 = ~n11511 ;
  assign n12151 = n29496 & n11652 ;
  assign n12152 = n12150 & n12151 ;
  assign n12291 = n12150 | n12151 ;
  assign n29497 = ~n12152 ;
  assign n12292 = n29497 & n12291 ;
  assign n12293 = n12290 & n12292 ;
  assign n12474 = n12290 | n12292 ;
  assign n29498 = ~n12293 ;
  assign n12475 = n29498 & n12474 ;
  assign n12873 = n12304 | n12872 ;
  assign n29499 = ~n12873 ;
  assign n12874 = n12475 & n29499 ;
  assign n29500 = ~n12475 ;
  assign n13161 = n29500 & n12873 ;
  assign n13162 = n12874 | n13161 ;
  assign n13163 = n13160 & n13162 ;
  assign n13396 = n13160 | n13162 ;
  assign n29501 = ~n13163 ;
  assign n13397 = n29501 & n13396 ;
  assign n13398 = n13395 & n13397 ;
  assign n13894 = n13395 | n13397 ;
  assign n29502 = ~n13398 ;
  assign n13895 = n29502 & n13894 ;
  assign n29503 = ~n13893 ;
  assign n13897 = n29503 & n13895 ;
  assign n29504 = ~n13895 ;
  assign n13898 = n13893 & n29504 ;
  assign n13899 = n13897 | n13898 ;
  assign n13909 = n13900 & n13907 ;
  assign n14177 = n13924 & n14176 ;
  assign n14178 = n13925 | n14177 ;
  assign n14179 = n13914 & n14178 ;
  assign n14180 = n13909 | n14179 ;
  assign n14181 = n13899 | n14180 ;
  assign n14182 = n13899 & n14180 ;
  assign n29505 = ~n14182 ;
  assign n14790 = n14181 & n29505 ;
  assign n5315 = n1522 & n5302 ;
  assign n5280 = x[85] & n5240 ;
  assign n6238 = x[86] & n6179 ;
  assign n14791 = n5280 | n6238 ;
  assign n14792 = x[87] & n5238 ;
  assign n14793 = n14791 | n14792 ;
  assign n14794 = n5315 | n14793 ;
  assign n29506 = ~n14794 ;
  assign n14795 = x[23] & n29506 ;
  assign n14796 = n28221 & n14794 ;
  assign n14797 = n14795 | n14796 ;
  assign n14798 = n14790 & n14797 ;
  assign n13896 = n13893 & n13895 ;
  assign n14693 = n13893 | n13895 ;
  assign n29507 = ~n13896 ;
  assign n14694 = n29507 & n14693 ;
  assign n29508 = ~n14180 ;
  assign n14695 = n29508 & n14694 ;
  assign n29509 = ~n14694 ;
  assign n15720 = n14180 & n29509 ;
  assign n15721 = n14695 | n15720 ;
  assign n15722 = n14797 | n15721 ;
  assign n29510 = ~n14798 ;
  assign n15801 = n29510 & n15722 ;
  assign n29511 = ~n15801 ;
  assign n15802 = n15116 & n29511 ;
  assign n15723 = n14797 & n15721 ;
  assign n15724 = n14807 & n14810 ;
  assign n15796 = n14823 | n15795 ;
  assign n15797 = n15725 & n15796 ;
  assign n15798 = n15724 | n15797 ;
  assign n15799 = n15722 & n15798 ;
  assign n15800 = n15723 | n15799 ;
  assign n29512 = ~n15800 ;
  assign n15803 = n15722 & n29512 ;
  assign n15804 = n15802 | n15803 ;
  assign n7202 = n1482 & n7162 ;
  assign n7114 = x[88] & n7100 ;
  assign n7676 = x[89] & n7647 ;
  assign n15805 = n7114 | n7676 ;
  assign n15806 = x[90] & n7098 ;
  assign n15807 = n15805 | n15806 ;
  assign n15808 = n7202 | n15807 ;
  assign n29513 = ~n15808 ;
  assign n15809 = x[20] & n29513 ;
  assign n15810 = n28114 & n15808 ;
  assign n15811 = n15809 | n15810 ;
  assign n29514 = ~n15811 ;
  assign n15812 = n15804 & n29514 ;
  assign n29515 = ~n15804 ;
  assign n16484 = n29515 & n15811 ;
  assign n16485 = n15812 | n16484 ;
  assign n16486 = n16483 & n16485 ;
  assign n16727 = n16483 | n16485 ;
  assign n29516 = ~n16486 ;
  assign n16728 = n29516 & n16727 ;
  assign n16729 = n16726 & n16728 ;
  assign n17145 = n16726 | n16728 ;
  assign n29517 = ~n16729 ;
  assign n17146 = n29517 & n17145 ;
  assign n17147 = n17144 & n17146 ;
  assign n17695 = n17144 | n17146 ;
  assign n29518 = ~n17147 ;
  assign n17696 = n29518 & n17695 ;
  assign n17697 = n17694 & n17696 ;
  assign n18223 = n17694 | n17696 ;
  assign n29519 = ~n17697 ;
  assign n18739 = n29519 & n18223 ;
  assign n29520 = ~n18222 ;
  assign n18741 = n29520 & n18739 ;
  assign n29521 = ~n18739 ;
  assign n18938 = n18222 & n29521 ;
  assign n18939 = n18741 | n18938 ;
  assign n29522 = ~n18937 ;
  assign n18941 = n29522 & n18939 ;
  assign n29523 = ~n18939 ;
  assign n18942 = n18937 & n29523 ;
  assign n18943 = n18941 | n18942 ;
  assign n19515 = n18966 | n19514 ;
  assign n19516 = n18956 & n19515 ;
  assign n19517 = n18953 | n19516 ;
  assign n19518 = n18943 | n19517 ;
  assign n19519 = n18943 & n19517 ;
  assign n29524 = ~n19519 ;
  assign n20861 = n19518 & n29524 ;
  assign n29525 = ~n20223 ;
  assign n20862 = n29525 & n20861 ;
  assign n29526 = ~n20861 ;
  assign n20863 = n20223 & n29526 ;
  assign n20864 = n20862 | n20863 ;
  assign n21270 = n20233 | n21119 ;
  assign n21271 = n21269 & n21270 ;
  assign n21272 = n21120 | n21271 ;
  assign n29527 = ~n20864 ;
  assign n21273 = n29527 & n21272 ;
  assign n29528 = ~n21272 ;
  assign n21383 = n20864 & n29528 ;
  assign n21384 = n21273 | n21383 ;
  assign n29529 = ~n21382 ;
  assign n21987 = n29529 & n21384 ;
  assign n29530 = ~n21384 ;
  assign n22273 = n21382 & n29530 ;
  assign n22274 = n21987 | n22273 ;
  assign n22275 = n22272 | n22274 ;
  assign n22276 = n22272 & n22274 ;
  assign n29531 = ~n22276 ;
  assign n23019 = n22275 & n29531 ;
  assign n585 = n583 & n584 ;
  assign n586 = n27620 | n585 ;
  assign n24903 = x[107] & x[108] ;
  assign n587 = x[107] | x[108] ;
  assign n29532 = ~n24903 ;
  assign n3873 = n29532 & n587 ;
  assign n3874 = n586 & n3873 ;
  assign n3875 = n586 | n3873 ;
  assign n29533 = ~n3874 ;
  assign n3876 = n29533 & n3875 ;
  assign n19710 = n3876 & n19656 ;
  assign n19736 = x[106] & n19723 ;
  assign n19891 = x[107] & n19829 ;
  assign n23020 = n19736 | n19891 ;
  assign n23021 = x[108] & n19655 ;
  assign n23022 = n23020 | n23021 ;
  assign n23023 = n19710 | n23022 ;
  assign n29534 = ~n23023 ;
  assign n23024 = x[2] & n29534 ;
  assign n23025 = n27790 & n23023 ;
  assign n23026 = n23024 | n23025 ;
  assign n23027 = n23019 | n23026 ;
  assign n23028 = n23019 & n23026 ;
  assign n29535 = ~n23028 ;
  assign n23029 = n23027 & n29535 ;
  assign n23030 = n23018 & n23029 ;
  assign n27687 = n23018 | n23029 ;
  assign n29536 = ~n23030 ;
  assign n173 = n29536 & n27687 ;
  assign n23031 = n23028 | n23030 ;
  assign n21385 = n21382 & n21384 ;
  assign n21975 = n21972 & n21974 ;
  assign n21976 = n21416 | n21975 ;
  assign n21979 = n21403 & n21978 ;
  assign n21981 = n21403 | n21978 ;
  assign n29537 = ~n21979 ;
  assign n21982 = n29537 & n21981 ;
  assign n21983 = n21976 & n21982 ;
  assign n21984 = n21406 | n21983 ;
  assign n21985 = n21395 & n21984 ;
  assign n21986 = n21396 | n21985 ;
  assign n21988 = n21382 | n21384 ;
  assign n29538 = ~n21385 ;
  assign n21989 = n29538 & n21988 ;
  assign n21990 = n21986 & n21989 ;
  assign n21991 = n21385 | n21990 ;
  assign n18940 = n18937 & n18939 ;
  assign n19520 = n18940 | n19519 ;
  assign n12751 = n2466 & n12695 ;
  assign n12659 = x[98] & n12633 ;
  assign n14388 = x[99] & n13533 ;
  assign n18923 = n12659 | n14388 ;
  assign n18924 = x[100] & n12631 ;
  assign n18925 = n18923 | n18924 ;
  assign n18926 = n12751 | n18925 ;
  assign n29539 = ~n18926 ;
  assign n18927 = x[11] & n29539 ;
  assign n18928 = n27892 & n18926 ;
  assign n18929 = n18927 | n18928 ;
  assign n18224 = n18222 & n18223 ;
  assign n18225 = n17697 | n18224 ;
  assign n10575 = n2438 & n10542 ;
  assign n10512 = x[95] & n10481 ;
  assign n11870 = x[96] & n11232 ;
  assign n17678 = n10512 | n11870 ;
  assign n17679 = x[97] & n10479 ;
  assign n17680 = n17678 | n17679 ;
  assign n17681 = n10575 | n17680 ;
  assign n29540 = ~n17681 ;
  assign n17682 = x[14] & n29540 ;
  assign n17683 = n27956 & n17681 ;
  assign n17684 = n17682 | n17683 ;
  assign n17148 = n16729 | n17147 ;
  assign n15813 = n15804 & n15811 ;
  assign n16487 = n15813 | n16486 ;
  assign n7197 = n2046 & n7162 ;
  assign n7145 = x[89] & n7100 ;
  assign n7688 = x[90] & n7647 ;
  assign n15710 = n7145 | n7688 ;
  assign n15711 = x[91] & n7098 ;
  assign n15712 = n15710 | n15711 ;
  assign n15713 = n7197 | n15712 ;
  assign n29541 = ~n15713 ;
  assign n15714 = x[20] & n29541 ;
  assign n15715 = n28114 & n15713 ;
  assign n15716 = n15714 | n15715 ;
  assign n15117 = n14790 | n14797 ;
  assign n15118 = n15116 & n15117 ;
  assign n15119 = n14798 | n15118 ;
  assign n1242 = n452 & n1239 ;
  assign n346 = x[83] & n330 ;
  assign n438 = x[84] & n390 ;
  assign n13874 = n346 | n438 ;
  assign n13875 = x[85] & n322 ;
  assign n13876 = n13874 | n13875 ;
  assign n13877 = n1242 | n13876 ;
  assign n29542 = ~n13877 ;
  assign n13878 = x[26] & n29542 ;
  assign n13879 = n28342 & n13877 ;
  assign n13880 = n13878 | n13879 ;
  assign n13399 = n13163 | n13398 ;
  assign n12144 = n11510 & n11651 ;
  assign n12153 = n12144 | n12152 ;
  assign n4050 = n2750 & n4041 ;
  assign n3923 = x[74] & n3910 ;
  assign n3987 = x[75] & n3975 ;
  assign n11492 = n3923 | n3987 ;
  assign n11493 = x[76] & n3906 ;
  assign n11494 = n11492 | n11493 ;
  assign n11495 = n4050 | n11494 ;
  assign n29543 = ~n11495 ;
  assign n11496 = x[35] & n29543 ;
  assign n11497 = n28822 & n11495 ;
  assign n11498 = n11496 | n11497 ;
  assign n10945 = n10941 & n10943 ;
  assign n11045 = n10945 | n11044 ;
  assign n5981 = n3162 & n5976 ;
  assign n3043 = x[68] & n3031 ;
  assign n3115 = x[69] & n3096 ;
  assign n10206 = n3043 | n3115 ;
  assign n10207 = x[70] & n3027 ;
  assign n10208 = n10206 | n10207 ;
  assign n10209 = n5981 | n10208 ;
  assign n29544 = ~n10209 ;
  assign n10210 = x[41] & n29544 ;
  assign n10211 = n29184 & n10209 ;
  assign n10212 = n10210 | n10211 ;
  assign n27700 = x[44] & x[45] ;
  assign n2171 = x[44] | x[45] ;
  assign n29545 = ~n27700 ;
  assign n2172 = n29545 & n2171 ;
  assign n9026 = x[64] & n2172 ;
  assign n9576 = n9567 & n9574 ;
  assign n9577 = n9026 & n9576 ;
  assign n9578 = n9026 | n9576 ;
  assign n29546 = ~n9577 ;
  assign n9579 = n29546 & n9578 ;
  assign n6497 = n2635 & n6494 ;
  assign n2550 = x[65] & n2492 ;
  assign n2567 = x[66] & n2557 ;
  assign n9580 = n2550 | n2567 ;
  assign n9581 = x[67] & n2488 ;
  assign n9582 = n9580 | n9581 ;
  assign n9583 = n6497 | n9582 ;
  assign n29547 = ~n9583 ;
  assign n9584 = x[44] & n29547 ;
  assign n9585 = n29400 & n9583 ;
  assign n9586 = n9584 | n9585 ;
  assign n29548 = ~n9586 ;
  assign n9587 = n9579 & n29548 ;
  assign n29549 = ~n9579 ;
  assign n10213 = n29549 & n9586 ;
  assign n10214 = n9587 | n10213 ;
  assign n10215 = n10212 & n10214 ;
  assign n10216 = n10212 | n10214 ;
  assign n29550 = ~n10215 ;
  assign n10217 = n29550 & n10216 ;
  assign n10228 = n10219 & n10226 ;
  assign n10280 = n10276 & n10278 ;
  assign n10281 = n10228 | n10280 ;
  assign n29551 = ~n10281 ;
  assign n10282 = n10217 & n29551 ;
  assign n29552 = ~n10217 ;
  assign n10925 = n29552 & n10281 ;
  assign n10926 = n10282 | n10925 ;
  assign n3736 = n3574 & n3733 ;
  assign n3452 = x[71] & n3443 ;
  assign n3541 = x[72] & n3508 ;
  assign n10927 = n3452 | n3541 ;
  assign n10928 = x[73] & n3439 ;
  assign n10929 = n10927 | n10928 ;
  assign n10930 = n3736 | n10929 ;
  assign n29553 = ~n10930 ;
  assign n10931 = x[38] & n29553 ;
  assign n10932 = n28996 & n10930 ;
  assign n10933 = n10931 | n10932 ;
  assign n10934 = n10926 & n10933 ;
  assign n11046 = n10926 | n10933 ;
  assign n29554 = ~n10934 ;
  assign n11047 = n29554 & n11046 ;
  assign n11048 = n11045 & n11047 ;
  assign n11499 = n11045 | n11047 ;
  assign n29555 = ~n11048 ;
  assign n11500 = n29555 & n11499 ;
  assign n29556 = ~n11498 ;
  assign n11655 = n29556 & n11500 ;
  assign n29557 = ~n11500 ;
  assign n12154 = n11498 & n29557 ;
  assign n12155 = n11655 | n12154 ;
  assign n12156 = n12153 | n12155 ;
  assign n12157 = n12153 & n12155 ;
  assign n29558 = ~n12157 ;
  assign n12274 = n12156 & n29558 ;
  assign n1743 = n779 & n1741 ;
  assign n711 = x[77] & n663 ;
  assign n744 = x[78] & n720 ;
  assign n12275 = n711 | n744 ;
  assign n12276 = x[79] & n652 ;
  assign n12277 = n12275 | n12276 ;
  assign n12278 = n1743 | n12277 ;
  assign n29559 = ~n12278 ;
  assign n12279 = x[32] & n29559 ;
  assign n12280 = n28658 & n12278 ;
  assign n12281 = n12279 | n12280 ;
  assign n29560 = ~n12281 ;
  assign n12478 = n12274 & n29560 ;
  assign n29561 = ~n12274 ;
  assign n12479 = n29561 & n12281 ;
  assign n12480 = n12478 | n12479 ;
  assign n12875 = n12474 & n12873 ;
  assign n12876 = n12293 | n12875 ;
  assign n29562 = ~n12480 ;
  assign n12877 = n29562 & n12876 ;
  assign n29563 = ~n12876 ;
  assign n13143 = n12480 & n29563 ;
  assign n13144 = n12877 | n13143 ;
  assign n4639 = n1003 & n4632 ;
  assign n4559 = x[80] & n4514 ;
  assign n4618 = x[81] & n4572 ;
  assign n13145 = n4559 | n4618 ;
  assign n13146 = x[82] & n4504 ;
  assign n13147 = n13145 | n13146 ;
  assign n13148 = n4639 | n13147 ;
  assign n29564 = ~n13148 ;
  assign n13149 = x[29] & n29564 ;
  assign n13150 = n28483 & n13148 ;
  assign n13151 = n13149 | n13150 ;
  assign n13152 = n13144 | n13151 ;
  assign n13153 = n13144 & n13151 ;
  assign n29565 = ~n13153 ;
  assign n13794 = n13152 & n29565 ;
  assign n29566 = ~n13399 ;
  assign n13796 = n29566 & n13794 ;
  assign n29567 = ~n13794 ;
  assign n13881 = n13399 & n29567 ;
  assign n13882 = n13796 | n13881 ;
  assign n13883 = n13880 & n13882 ;
  assign n13885 = n13880 | n13882 ;
  assign n29568 = ~n13883 ;
  assign n13886 = n29568 & n13885 ;
  assign n14741 = n13913 | n14740 ;
  assign n14742 = n14694 & n14741 ;
  assign n14743 = n13896 | n14742 ;
  assign n29569 = ~n14743 ;
  assign n14744 = n13886 & n29569 ;
  assign n29570 = ~n13886 ;
  assign n14779 = n29570 & n14743 ;
  assign n14780 = n14744 | n14779 ;
  assign n5316 = n1720 & n5302 ;
  assign n5253 = x[86] & n5240 ;
  assign n6240 = x[87] & n6179 ;
  assign n14781 = n5253 | n6240 ;
  assign n14782 = x[88] & n5238 ;
  assign n14783 = n14781 | n14782 ;
  assign n14784 = n5316 | n14783 ;
  assign n29571 = ~n14784 ;
  assign n14785 = x[23] & n29571 ;
  assign n14786 = n28221 & n14784 ;
  assign n14787 = n14785 | n14786 ;
  assign n14788 = n14780 | n14787 ;
  assign n14789 = n14780 & n14787 ;
  assign n29572 = ~n14789 ;
  assign n15120 = n14788 & n29572 ;
  assign n29573 = ~n15119 ;
  assign n15121 = n29573 & n15120 ;
  assign n29574 = ~n15120 ;
  assign n15717 = n15119 & n29574 ;
  assign n15718 = n15121 | n15717 ;
  assign n29575 = ~n15716 ;
  assign n16182 = n29575 & n15718 ;
  assign n29576 = ~n15718 ;
  assign n16488 = n15716 & n29576 ;
  assign n16489 = n16182 | n16488 ;
  assign n16490 = n16487 | n16489 ;
  assign n16491 = n16487 & n16489 ;
  assign n29577 = ~n16491 ;
  assign n16711 = n16490 & n29577 ;
  assign n8740 = n2410 & n8706 ;
  assign n8663 = x[92] & n8645 ;
  assign n9880 = x[93] & n9278 ;
  assign n16712 = n8663 | n9880 ;
  assign n16713 = x[94] & n8643 ;
  assign n16714 = n16712 | n16713 ;
  assign n16715 = n8740 | n16714 ;
  assign n29578 = ~n16715 ;
  assign n16716 = x[17] & n29578 ;
  assign n16717 = n28039 & n16715 ;
  assign n16718 = n16716 | n16717 ;
  assign n16719 = n16711 & n16718 ;
  assign n17149 = n16711 | n16718 ;
  assign n29579 = ~n16719 ;
  assign n17476 = n29579 & n17149 ;
  assign n29580 = ~n17148 ;
  assign n17478 = n29580 & n17476 ;
  assign n29581 = ~n17476 ;
  assign n17685 = n17148 & n29581 ;
  assign n17686 = n17478 | n17685 ;
  assign n29582 = ~n17684 ;
  assign n18226 = n29582 & n17686 ;
  assign n29583 = ~n17686 ;
  assign n18743 = n17684 & n29583 ;
  assign n18744 = n18226 | n18743 ;
  assign n29584 = ~n18744 ;
  assign n18746 = n18225 & n29584 ;
  assign n29585 = ~n18225 ;
  assign n19521 = n29585 & n18744 ;
  assign n19522 = n18746 | n19521 ;
  assign n19523 = n18929 & n19522 ;
  assign n18737 = n18219 & n18735 ;
  assign n18738 = n17707 | n18737 ;
  assign n18740 = n18738 & n18739 ;
  assign n18742 = n17697 | n18740 ;
  assign n18745 = n18742 | n18744 ;
  assign n18747 = n18742 & n18744 ;
  assign n29586 = ~n18747 ;
  assign n18922 = n18745 & n29586 ;
  assign n19524 = n18922 | n18929 ;
  assign n29587 = ~n19523 ;
  assign n19525 = n29587 & n19524 ;
  assign n19526 = n19520 & n19525 ;
  assign n20202 = n19520 | n19525 ;
  assign n29588 = ~n19526 ;
  assign n20203 = n29588 & n20202 ;
  assign n15351 = n2626 & n15308 ;
  assign n15293 = x[101] & n15246 ;
  assign n17323 = x[102] & n16288 ;
  assign n20204 = n15293 | n17323 ;
  assign n20205 = x[103] & n15244 ;
  assign n20206 = n20204 | n20205 ;
  assign n20207 = n15351 | n20206 ;
  assign n29589 = ~n20207 ;
  assign n20208 = x[8] & n29589 ;
  assign n20209 = n27845 & n20207 ;
  assign n20210 = n20208 | n20209 ;
  assign n20212 = n20203 & n20210 ;
  assign n20213 = n20203 | n20210 ;
  assign n29590 = ~n20212 ;
  assign n20214 = n29590 & n20213 ;
  assign n21117 = n20223 & n20861 ;
  assign n20055 = n18937 | n18939 ;
  assign n29591 = ~n18940 ;
  assign n20056 = n29591 & n20055 ;
  assign n29592 = ~n19517 ;
  assign n20057 = n29592 & n20056 ;
  assign n29593 = ~n20056 ;
  assign n20215 = n19517 & n29593 ;
  assign n20216 = n20057 | n20215 ;
  assign n20224 = n20216 | n20223 ;
  assign n20225 = n20216 & n20223 ;
  assign n29594 = ~n20225 ;
  assign n21274 = n20224 & n29594 ;
  assign n21275 = n21272 & n21274 ;
  assign n21276 = n21117 | n21275 ;
  assign n29595 = ~n21276 ;
  assign n21277 = n20214 & n29595 ;
  assign n29596 = ~n20214 ;
  assign n21361 = n29596 & n21276 ;
  assign n21362 = n21277 | n21361 ;
  assign n18437 = n3223 & n18392 ;
  assign n18361 = x[104] & n18329 ;
  assign n18551 = x[105] & n18514 ;
  assign n21363 = n18361 | n18551 ;
  assign n21364 = x[106] & n18327 ;
  assign n21365 = n21363 | n21364 ;
  assign n21366 = n18437 | n21365 ;
  assign n29597 = ~n21366 ;
  assign n21367 = x[5] & n29597 ;
  assign n21368 = n27813 & n21366 ;
  assign n21369 = n21367 | n21368 ;
  assign n21370 = n21362 | n21369 ;
  assign n21371 = n21362 & n21369 ;
  assign n29598 = ~n21371 ;
  assign n22100 = n21370 & n29598 ;
  assign n29599 = ~n21991 ;
  assign n22101 = n29599 & n22100 ;
  assign n29600 = ~n22100 ;
  assign n22380 = n21991 & n29600 ;
  assign n22381 = n22101 | n22380 ;
  assign n588 = n586 & n587 ;
  assign n589 = n24903 | n588 ;
  assign n27619 = x[108] & x[109] ;
  assign n590 = x[108] | x[109] ;
  assign n29601 = ~n27619 ;
  assign n3636 = n29601 & n590 ;
  assign n3637 = n589 | n3636 ;
  assign n3638 = n589 & n3636 ;
  assign n29602 = ~n3638 ;
  assign n3639 = n3637 & n29602 ;
  assign n19664 = n3639 & n19656 ;
  assign n19778 = x[107] & n19723 ;
  assign n19868 = x[108] & n19829 ;
  assign n22382 = n19778 | n19868 ;
  assign n22383 = x[109] & n19655 ;
  assign n22384 = n22382 | n22383 ;
  assign n22385 = n19664 | n22384 ;
  assign n29603 = ~n22385 ;
  assign n22386 = x[2] & n29603 ;
  assign n22387 = n27790 & n22385 ;
  assign n22388 = n22386 | n22387 ;
  assign n22389 = n22381 | n22388 ;
  assign n22390 = n22381 & n22388 ;
  assign n29604 = ~n22390 ;
  assign n23032 = n22389 & n29604 ;
  assign n23033 = n23031 | n23032 ;
  assign n23034 = n23031 & n23032 ;
  assign n29605 = ~n23034 ;
  assign n174 = n23033 & n29605 ;
  assign n29606 = ~n20210 ;
  assign n20211 = n20203 & n29606 ;
  assign n29607 = ~n20203 ;
  assign n21115 = n29607 & n20210 ;
  assign n21116 = n20211 | n21115 ;
  assign n21279 = n21116 & n21276 ;
  assign n21280 = n20212 | n21279 ;
  assign n18930 = n18922 & n18929 ;
  assign n19527 = n18930 | n19526 ;
  assign n17687 = n17684 & n17686 ;
  assign n18227 = n17684 | n17686 ;
  assign n29608 = ~n17687 ;
  assign n18228 = n29608 & n18227 ;
  assign n18229 = n18225 & n18228 ;
  assign n18230 = n17687 | n18229 ;
  assign n10567 = n2841 & n10542 ;
  assign n10498 = x[96] & n10481 ;
  assign n11871 = x[97] & n11232 ;
  assign n17665 = n10498 | n11871 ;
  assign n17666 = x[98] & n10479 ;
  assign n17667 = n17665 | n17666 ;
  assign n17668 = n10567 | n17667 ;
  assign n29609 = ~n17668 ;
  assign n17669 = x[14] & n29609 ;
  assign n17670 = n27956 & n17668 ;
  assign n17671 = n17669 | n17670 ;
  assign n7177 = n1841 & n7162 ;
  assign n7153 = x[90] & n7100 ;
  assign n7710 = x[91] & n7647 ;
  assign n15700 = n7153 | n7710 ;
  assign n15701 = x[92] & n7098 ;
  assign n15702 = n15700 | n15701 ;
  assign n15703 = n7177 | n15702 ;
  assign n29610 = ~n15703 ;
  assign n15704 = x[20] & n29610 ;
  assign n15705 = n28114 & n15703 ;
  assign n15706 = n15704 | n15705 ;
  assign n15122 = n15119 & n15120 ;
  assign n15123 = n14789 | n15122 ;
  assign n1216 = n452 & n1213 ;
  assign n347 = x[84] & n330 ;
  assign n436 = x[85] & n390 ;
  assign n13861 = n347 | n436 ;
  assign n13862 = x[86] & n322 ;
  assign n13863 = n13861 | n13862 ;
  assign n13864 = n1216 | n13863 ;
  assign n29611 = ~n13864 ;
  assign n13865 = x[26] & n29611 ;
  assign n13866 = n28342 & n13864 ;
  assign n13867 = n13865 | n13866 ;
  assign n1271 = n779 & n1270 ;
  assign n693 = x[78] & n663 ;
  assign n763 = x[79] & n720 ;
  assign n12261 = n693 | n763 ;
  assign n12262 = x[80] & n652 ;
  assign n12263 = n12261 | n12262 ;
  assign n12264 = n1271 | n12263 ;
  assign n29612 = ~n12264 ;
  assign n12265 = x[32] & n29612 ;
  assign n12266 = n28658 & n12264 ;
  assign n12267 = n12265 | n12266 ;
  assign n11501 = n11498 & n11500 ;
  assign n12158 = n11501 | n12157 ;
  assign n4795 = n3162 & n4790 ;
  assign n3045 = x[69] & n3031 ;
  assign n3151 = x[70] & n3096 ;
  assign n10193 = n3045 | n3151 ;
  assign n10194 = x[71] & n3027 ;
  assign n10195 = n10193 | n10194 ;
  assign n10196 = n4795 | n10195 ;
  assign n29613 = ~n10196 ;
  assign n10197 = x[41] & n29613 ;
  assign n10198 = n29184 & n10196 ;
  assign n10199 = n10197 | n10198 ;
  assign n9588 = n9579 & n9586 ;
  assign n9589 = n9577 | n9588 ;
  assign n6414 = n2635 & n6408 ;
  assign n2501 = x[66] & n2492 ;
  assign n2570 = x[67] & n2557 ;
  assign n9547 = n2501 | n2570 ;
  assign n9548 = x[68] & n2488 ;
  assign n9549 = n9547 | n9548 ;
  assign n9550 = n6414 | n9549 ;
  assign n9551 = x[44] | n9550 ;
  assign n9552 = x[44] & n9550 ;
  assign n29614 = ~n9552 ;
  assign n9553 = n9551 & n29614 ;
  assign n29615 = ~n9026 ;
  assign n9027 = x[47] & n29615 ;
  assign n27701 = x[46] & x[47] ;
  assign n2173 = x[46] | x[47] ;
  assign n29616 = ~n27701 ;
  assign n2174 = n29616 & n2173 ;
  assign n2321 = n2172 & n2174 ;
  assign n6442 = n2321 & n6437 ;
  assign n29617 = ~n2174 ;
  assign n2175 = n2172 & n29617 ;
  assign n9028 = x[65] & n2175 ;
  assign n27703 = x[45] & x[46] ;
  assign n2176 = x[45] | x[46] ;
  assign n29618 = ~n27703 ;
  assign n2177 = n29618 & n2176 ;
  assign n29619 = ~n2172 ;
  assign n2244 = n29619 & n2177 ;
  assign n9029 = x[64] & n2244 ;
  assign n9030 = n9028 | n9029 ;
  assign n9031 = n6442 | n9030 ;
  assign n29620 = ~n9031 ;
  assign n9032 = x[47] & n29620 ;
  assign n29621 = ~x[47] ;
  assign n9033 = n29621 & n9031 ;
  assign n9034 = n9032 | n9033 ;
  assign n29622 = ~n9034 ;
  assign n9035 = n9027 & n29622 ;
  assign n29623 = ~n9027 ;
  assign n9554 = n29623 & n9034 ;
  assign n9555 = n9035 | n9554 ;
  assign n9556 = n9553 & n9555 ;
  assign n9590 = n9553 | n9555 ;
  assign n29624 = ~n9556 ;
  assign n9591 = n29624 & n9590 ;
  assign n29625 = ~n9589 ;
  assign n9592 = n29625 & n9591 ;
  assign n29626 = ~n9591 ;
  assign n10200 = n9589 & n29626 ;
  assign n10201 = n9592 | n10200 ;
  assign n29627 = ~n10199 ;
  assign n10202 = n29627 & n10201 ;
  assign n29628 = ~n10201 ;
  assign n10204 = n10199 & n29628 ;
  assign n10205 = n10202 | n10204 ;
  assign n10283 = n10217 & n10281 ;
  assign n10284 = n10215 | n10283 ;
  assign n29629 = ~n10284 ;
  assign n10285 = n10205 & n29629 ;
  assign n29630 = ~n10205 ;
  assign n10915 = n29630 & n10284 ;
  assign n10916 = n10285 | n10915 ;
  assign n3583 = n2722 & n3574 ;
  assign n3459 = x[72] & n3443 ;
  assign n3522 = x[73] & n3508 ;
  assign n10917 = n3459 | n3522 ;
  assign n10918 = x[74] & n3439 ;
  assign n10919 = n10917 | n10918 ;
  assign n10920 = n3583 | n10919 ;
  assign n29631 = ~n10920 ;
  assign n10921 = x[38] & n29631 ;
  assign n10922 = n28996 & n10920 ;
  assign n10923 = n10921 | n10922 ;
  assign n11050 = n10916 | n10923 ;
  assign n10924 = n10916 & n10923 ;
  assign n11476 = n11045 & n11046 ;
  assign n11477 = n10934 | n11476 ;
  assign n11478 = n11050 & n11477 ;
  assign n11479 = n10924 | n11478 ;
  assign n29632 = ~n11479 ;
  assign n11480 = n11050 & n29632 ;
  assign n11049 = n10934 | n11048 ;
  assign n29633 = ~n10924 ;
  assign n11051 = n29633 & n11050 ;
  assign n29634 = ~n11051 ;
  assign n11481 = n11049 & n29634 ;
  assign n11482 = n11480 | n11481 ;
  assign n4047 = n1775 & n4041 ;
  assign n3926 = x[75] & n3910 ;
  assign n3988 = x[76] & n3975 ;
  assign n11483 = n3926 | n3988 ;
  assign n11484 = x[77] & n3906 ;
  assign n11485 = n11483 | n11484 ;
  assign n11486 = n4047 | n11485 ;
  assign n29635 = ~n11486 ;
  assign n11487 = x[35] & n29635 ;
  assign n11488 = n28822 & n11486 ;
  assign n11489 = n11487 | n11488 ;
  assign n11490 = n11482 | n11489 ;
  assign n11491 = n11482 & n11489 ;
  assign n29636 = ~n11491 ;
  assign n12159 = n11490 & n29636 ;
  assign n12160 = n12158 & n12159 ;
  assign n12268 = n12158 | n12159 ;
  assign n29637 = ~n12160 ;
  assign n12269 = n29637 & n12268 ;
  assign n29638 = ~n12267 ;
  assign n12271 = n29638 & n12269 ;
  assign n29639 = ~n12269 ;
  assign n12863 = n12267 & n29639 ;
  assign n12864 = n12271 | n12863 ;
  assign n12283 = n12274 & n12281 ;
  assign n12282 = n12274 | n12281 ;
  assign n29640 = ~n12283 ;
  assign n12878 = n12282 & n29640 ;
  assign n12879 = n12876 & n12878 ;
  assign n12880 = n12283 | n12879 ;
  assign n12881 = n12864 | n12880 ;
  assign n12883 = n12864 & n12880 ;
  assign n29641 = ~n12883 ;
  assign n13128 = n12881 & n29641 ;
  assign n4640 = n1057 & n4632 ;
  assign n4558 = x[81] & n4514 ;
  assign n4597 = x[82] & n4572 ;
  assign n13129 = n4558 | n4597 ;
  assign n13130 = x[83] & n4504 ;
  assign n13131 = n13129 | n13130 ;
  assign n13132 = n4640 | n13131 ;
  assign n29642 = ~n13132 ;
  assign n13133 = x[29] & n29642 ;
  assign n13134 = n28483 & n13132 ;
  assign n13135 = n13133 | n13134 ;
  assign n29643 = ~n13135 ;
  assign n13136 = n13128 & n29643 ;
  assign n29644 = ~n13128 ;
  assign n13761 = n29644 & n13135 ;
  assign n13762 = n13136 | n13761 ;
  assign n13775 = n13232 | n13774 ;
  assign n13776 = n13221 & n13775 ;
  assign n13777 = n13219 | n13776 ;
  assign n13778 = n13200 | n13207 ;
  assign n13779 = n13777 & n13778 ;
  assign n13780 = n13209 | n13779 ;
  assign n13782 = n13780 & n13781 ;
  assign n13784 = n13196 | n13782 ;
  assign n13788 = n13784 & n13786 ;
  assign n13789 = n13389 | n13788 ;
  assign n13790 = n13764 & n13789 ;
  assign n13791 = n13173 | n13790 ;
  assign n13792 = n13396 & n13791 ;
  assign n13793 = n13163 | n13792 ;
  assign n13795 = n13793 & n13794 ;
  assign n13797 = n13153 | n13795 ;
  assign n13799 = n13762 | n13797 ;
  assign n13800 = n13762 & n13797 ;
  assign n29645 = ~n13800 ;
  assign n13870 = n13799 & n29645 ;
  assign n29646 = ~n13867 ;
  assign n13871 = n29646 & n13870 ;
  assign n29647 = ~n13870 ;
  assign n13872 = n13867 & n29647 ;
  assign n13873 = n13871 | n13872 ;
  assign n14183 = n13896 | n14182 ;
  assign n14184 = n13886 & n14183 ;
  assign n14185 = n13883 | n14184 ;
  assign n14186 = n13873 | n14185 ;
  assign n14187 = n13873 & n14185 ;
  assign n29648 = ~n14187 ;
  assign n14764 = n14186 & n29648 ;
  assign n5318 = n1453 & n5302 ;
  assign n5278 = x[87] & n5240 ;
  assign n6266 = x[88] & n6179 ;
  assign n14765 = n5278 | n6266 ;
  assign n14766 = x[89] & n5238 ;
  assign n14767 = n14765 | n14766 ;
  assign n14768 = n5318 | n14767 ;
  assign n29649 = ~n14768 ;
  assign n14769 = x[23] & n29649 ;
  assign n14770 = n28221 & n14768 ;
  assign n14771 = n14769 | n14770 ;
  assign n29650 = ~n14771 ;
  assign n14772 = n14764 & n29650 ;
  assign n29651 = ~n14764 ;
  assign n15520 = n29651 & n14771 ;
  assign n15521 = n14772 | n15520 ;
  assign n15523 = n15123 | n15521 ;
  assign n15524 = n15123 & n15521 ;
  assign n29652 = ~n15524 ;
  assign n16187 = n15523 & n29652 ;
  assign n29653 = ~n15706 ;
  assign n16188 = n29653 & n16187 ;
  assign n29654 = ~n16187 ;
  assign n16190 = n15706 & n29654 ;
  assign n16191 = n16188 | n16190 ;
  assign n15719 = n15716 & n15718 ;
  assign n16492 = n15719 | n16491 ;
  assign n29655 = ~n16191 ;
  assign n16493 = n29655 & n16492 ;
  assign n29656 = ~n16492 ;
  assign n16701 = n16191 & n29656 ;
  assign n16702 = n16493 | n16701 ;
  assign n8742 = n2152 & n8706 ;
  assign n8665 = x[93] & n8645 ;
  assign n9879 = x[94] & n9278 ;
  assign n16703 = n8665 | n9879 ;
  assign n16704 = x[95] & n8643 ;
  assign n16705 = n16703 | n16704 ;
  assign n16706 = n8742 | n16705 ;
  assign n29657 = ~n16706 ;
  assign n16707 = x[17] & n29657 ;
  assign n16708 = n28039 & n16706 ;
  assign n16709 = n16707 | n16708 ;
  assign n16710 = n16702 & n16709 ;
  assign n17152 = n16702 | n16709 ;
  assign n29658 = ~n16710 ;
  assign n17153 = n29658 & n17152 ;
  assign n17140 = n16736 & n17138 ;
  assign n17470 = n16736 | n17138 ;
  assign n29659 = ~n17140 ;
  assign n17471 = n29659 & n17470 ;
  assign n17472 = n17468 & n17471 ;
  assign n17473 = n16739 | n17472 ;
  assign n17474 = n17145 & n17473 ;
  assign n17475 = n16729 | n17474 ;
  assign n17477 = n17475 & n17476 ;
  assign n17479 = n16719 | n17477 ;
  assign n29660 = ~n17479 ;
  assign n17480 = n17153 & n29660 ;
  assign n29661 = ~n17153 ;
  assign n17672 = n29661 & n17479 ;
  assign n17673 = n17480 | n17672 ;
  assign n17674 = n17671 & n17673 ;
  assign n18699 = n17671 | n17673 ;
  assign n29662 = ~n17674 ;
  assign n18700 = n29662 & n18699 ;
  assign n29663 = ~n18230 ;
  assign n18701 = n29663 & n18700 ;
  assign n29664 = ~n18700 ;
  assign n18907 = n18230 & n29664 ;
  assign n18908 = n18701 | n18907 ;
  assign n12722 = n2977 & n12695 ;
  assign n12675 = x[99] & n12633 ;
  assign n14402 = x[100] & n13533 ;
  assign n18909 = n12675 | n14402 ;
  assign n18910 = x[101] & n12631 ;
  assign n18911 = n18909 | n18910 ;
  assign n18912 = n12722 | n18911 ;
  assign n29665 = ~n18912 ;
  assign n18913 = x[11] & n29665 ;
  assign n18914 = n27892 & n18912 ;
  assign n18915 = n18913 | n18914 ;
  assign n18916 = n18908 | n18915 ;
  assign n18917 = n18908 & n18915 ;
  assign n29666 = ~n18917 ;
  assign n20053 = n18916 & n29666 ;
  assign n29667 = ~n19527 ;
  assign n20054 = n29667 & n20053 ;
  assign n29668 = ~n20053 ;
  assign n20192 = n19527 & n29668 ;
  assign n20193 = n20054 | n20192 ;
  assign n15330 = n3001 & n15308 ;
  assign n15299 = x[102] & n15246 ;
  assign n17305 = x[103] & n16288 ;
  assign n20194 = n15299 | n17305 ;
  assign n20195 = x[104] & n15244 ;
  assign n20196 = n20194 | n20195 ;
  assign n20197 = n15330 | n20196 ;
  assign n29669 = ~n20197 ;
  assign n20198 = x[8] & n29669 ;
  assign n20199 = n27845 & n20197 ;
  assign n20200 = n20198 | n20199 ;
  assign n20869 = n20193 | n20200 ;
  assign n29670 = ~n17671 ;
  assign n17675 = n29670 & n17673 ;
  assign n29671 = ~n17673 ;
  assign n17676 = n17671 & n29671 ;
  assign n17677 = n17675 | n17676 ;
  assign n18231 = n17677 | n18230 ;
  assign n18232 = n17677 & n18230 ;
  assign n29672 = ~n18232 ;
  assign n18918 = n18231 & n29672 ;
  assign n29673 = ~n18915 ;
  assign n18919 = n29673 & n18918 ;
  assign n29674 = ~n18918 ;
  assign n18920 = n18915 & n29674 ;
  assign n18921 = n18919 | n18920 ;
  assign n19528 = n18921 | n19527 ;
  assign n19529 = n18921 & n19527 ;
  assign n29675 = ~n19529 ;
  assign n21113 = n19528 & n29675 ;
  assign n21114 = n20200 & n21113 ;
  assign n29676 = ~n21114 ;
  assign n21346 = n20869 & n29676 ;
  assign n29677 = ~n21346 ;
  assign n21347 = n21280 & n29677 ;
  assign n20201 = n20193 & n20200 ;
  assign n20865 = n20859 & n20864 ;
  assign n20866 = n20225 | n20865 ;
  assign n20867 = n20214 & n20866 ;
  assign n20868 = n20212 | n20867 ;
  assign n20870 = n20868 & n20869 ;
  assign n20871 = n20201 | n20870 ;
  assign n29678 = ~n20871 ;
  assign n21348 = n20869 & n29678 ;
  assign n21349 = n21347 | n21348 ;
  assign n18451 = n3199 & n18392 ;
  assign n18368 = x[105] & n18329 ;
  assign n18569 = x[106] & n18514 ;
  assign n21350 = n18368 | n18569 ;
  assign n21351 = x[107] & n18327 ;
  assign n21352 = n21350 | n21351 ;
  assign n21353 = n18451 | n21352 ;
  assign n29679 = ~n21353 ;
  assign n21354 = x[5] & n29679 ;
  assign n21355 = n27813 & n21353 ;
  assign n21356 = n21354 | n21355 ;
  assign n29680 = ~n21356 ;
  assign n21357 = n21349 & n29680 ;
  assign n29681 = ~n21349 ;
  assign n21359 = n29681 & n21356 ;
  assign n21360 = n21357 | n21359 ;
  assign n21278 = n21116 | n21276 ;
  assign n29682 = ~n21279 ;
  assign n21372 = n21278 & n29682 ;
  assign n22099 = n21369 & n21372 ;
  assign n22277 = n21385 | n22276 ;
  assign n22278 = n22100 & n22277 ;
  assign n22279 = n22099 | n22278 ;
  assign n22280 = n21360 | n22279 ;
  assign n22281 = n21360 & n22279 ;
  assign n29683 = ~n22281 ;
  assign n22368 = n22280 & n29683 ;
  assign n591 = n589 & n590 ;
  assign n592 = n27619 | n591 ;
  assign n24735 = x[109] & x[110] ;
  assign n593 = x[109] | x[110] ;
  assign n29684 = ~n24735 ;
  assign n3612 = n29684 & n593 ;
  assign n3613 = n592 & n3612 ;
  assign n3614 = n592 | n3612 ;
  assign n29685 = ~n3613 ;
  assign n3615 = n29685 & n3614 ;
  assign n19704 = n3615 & n19656 ;
  assign n19734 = x[108] & n19723 ;
  assign n19883 = x[109] & n19829 ;
  assign n22369 = n19734 | n19883 ;
  assign n22370 = x[110] & n19655 ;
  assign n22371 = n22369 | n22370 ;
  assign n22372 = n19704 | n22371 ;
  assign n29686 = ~n22372 ;
  assign n22373 = x[2] & n29686 ;
  assign n22374 = n27790 & n22372 ;
  assign n22375 = n22373 | n22374 ;
  assign n29687 = ~n22375 ;
  assign n22376 = n22368 & n29687 ;
  assign n29688 = ~n22368 ;
  assign n22378 = n29688 & n22375 ;
  assign n22379 = n22376 | n22378 ;
  assign n23035 = n22390 | n23034 ;
  assign n23036 = n22379 & n23035 ;
  assign n27690 = n22379 | n23035 ;
  assign n29689 = ~n23036 ;
  assign n175 = n29689 & n27690 ;
  assign n594 = n592 & n593 ;
  assign n595 = n24735 | n594 ;
  assign n27618 = x[110] & x[111] ;
  assign n596 = x[110] | x[111] ;
  assign n29690 = ~n27618 ;
  assign n4243 = n29690 & n596 ;
  assign n29691 = ~n595 ;
  assign n4244 = n29691 & n4243 ;
  assign n29692 = ~n4243 ;
  assign n4245 = n595 & n29692 ;
  assign n4246 = n4244 | n4245 ;
  assign n19659 = n4246 & n19656 ;
  assign n19772 = x[109] & n19723 ;
  assign n19831 = x[110] & n19829 ;
  assign n22355 = n19772 | n19831 ;
  assign n22356 = x[111] & n19655 ;
  assign n22357 = n22355 | n22356 ;
  assign n22358 = n19659 | n22357 ;
  assign n29693 = ~n22358 ;
  assign n22359 = x[2] & n29693 ;
  assign n22360 = n27790 & n22358 ;
  assign n22361 = n22359 | n22360 ;
  assign n21358 = n21349 & n21356 ;
  assign n22282 = n21358 | n22281 ;
  assign n10555 = n2313 & n10542 ;
  assign n10509 = x[97] & n10481 ;
  assign n11899 = x[98] & n11232 ;
  assign n17652 = n10509 | n11899 ;
  assign n17653 = x[99] & n10479 ;
  assign n17654 = n17652 | n17653 ;
  assign n17655 = n10555 | n17654 ;
  assign n29694 = ~n17655 ;
  assign n17656 = x[14] & n29694 ;
  assign n17657 = n27956 & n17655 ;
  assign n17658 = n17656 | n17657 ;
  assign n17150 = n17148 & n17149 ;
  assign n17151 = n16719 | n17150 ;
  assign n17154 = n17151 & n17153 ;
  assign n17155 = n16710 | n17154 ;
  assign n8730 = n2000 & n8706 ;
  assign n8701 = x[94] & n8645 ;
  assign n9843 = x[95] & n9278 ;
  assign n16691 = n8701 | n9843 ;
  assign n16692 = x[96] & n8643 ;
  assign n16693 = n16691 | n16692 ;
  assign n16694 = n8730 | n16693 ;
  assign n29695 = ~n16694 ;
  assign n16695 = x[17] & n29695 ;
  assign n16696 = n28039 & n16694 ;
  assign n16697 = n16695 | n16696 ;
  assign n12270 = n12267 & n12269 ;
  assign n12272 = n12267 | n12269 ;
  assign n29696 = ~n12270 ;
  assign n12273 = n29696 & n12272 ;
  assign n29697 = ~n12880 ;
  assign n12882 = n12273 & n29697 ;
  assign n29698 = ~n12273 ;
  assign n13138 = n29698 & n12880 ;
  assign n13139 = n12882 | n13138 ;
  assign n13140 = n13135 | n13139 ;
  assign n13141 = n13135 & n13139 ;
  assign n29699 = ~n13141 ;
  assign n13142 = n13140 & n29699 ;
  assign n29700 = ~n13797 ;
  assign n13798 = n13142 & n29700 ;
  assign n29701 = ~n13142 ;
  assign n13859 = n29701 & n13797 ;
  assign n13860 = n13798 | n13859 ;
  assign n13868 = n13860 | n13867 ;
  assign n13869 = n13860 & n13867 ;
  assign n29702 = ~n13869 ;
  assign n14689 = n13868 & n29702 ;
  assign n29703 = ~n14185 ;
  assign n14690 = n29703 & n14689 ;
  assign n29704 = ~n14689 ;
  assign n14774 = n14185 & n29704 ;
  assign n14775 = n14690 | n14774 ;
  assign n14776 = n14771 | n14775 ;
  assign n14777 = n14771 & n14775 ;
  assign n29705 = ~n14777 ;
  assign n14778 = n14776 & n29705 ;
  assign n29706 = ~n15123 ;
  assign n15522 = n14778 & n29706 ;
  assign n29707 = ~n14778 ;
  assign n15707 = n29707 & n15123 ;
  assign n15708 = n15522 | n15707 ;
  assign n15709 = n15706 & n15708 ;
  assign n15823 = n15814 & n15821 ;
  assign n16175 = n16172 & n16174 ;
  assign n16176 = n15838 | n16175 ;
  assign n16177 = n15828 & n16176 ;
  assign n16178 = n15823 | n16177 ;
  assign n16179 = n15804 | n15811 ;
  assign n16180 = n16178 & n16179 ;
  assign n16181 = n15813 | n16180 ;
  assign n16183 = n15716 | n15718 ;
  assign n29708 = ~n15719 ;
  assign n16184 = n29708 & n16183 ;
  assign n16185 = n16181 & n16184 ;
  assign n16186 = n15719 | n16185 ;
  assign n16192 = n16186 & n16191 ;
  assign n16193 = n15709 | n16192 ;
  assign n7181 = n1685 & n7162 ;
  assign n7149 = x[91] & n7100 ;
  assign n7716 = x[92] & n7647 ;
  assign n15690 = n7149 | n7716 ;
  assign n15691 = x[93] & n7098 ;
  assign n15692 = n15690 | n15691 ;
  assign n15693 = n7181 | n15692 ;
  assign n29709 = ~n15693 ;
  assign n15694 = x[20] & n29709 ;
  assign n15695 = n28114 & n15693 ;
  assign n15696 = n15694 | n15695 ;
  assign n15525 = n14777 | n15524 ;
  assign n14188 = n13869 | n14187 ;
  assign n1031 = n779 & n1029 ;
  assign n676 = x[79] & n663 ;
  assign n762 = x[80] & n720 ;
  assign n12252 = n676 | n762 ;
  assign n12253 = x[81] & n652 ;
  assign n12254 = n12252 | n12253 ;
  assign n12255 = n1031 | n12254 ;
  assign n29710 = ~n12255 ;
  assign n12256 = x[32] & n29710 ;
  assign n12257 = n28658 & n12255 ;
  assign n12258 = n12256 | n12257 ;
  assign n12161 = n11491 | n12160 ;
  assign n4048 = n2084 & n4041 ;
  assign n3935 = x[76] & n3910 ;
  assign n3990 = x[77] & n3975 ;
  assign n11465 = n3935 | n3990 ;
  assign n11466 = x[78] & n3906 ;
  assign n11467 = n11465 | n11466 ;
  assign n11468 = n4048 | n11467 ;
  assign n29711 = ~n11468 ;
  assign n11469 = x[35] & n29711 ;
  assign n11470 = n28822 & n11468 ;
  assign n11471 = n11469 | n11470 ;
  assign n11052 = n11049 & n11050 ;
  assign n11053 = n10924 | n11052 ;
  assign n10203 = n10199 & n10201 ;
  assign n10286 = n10205 & n10284 ;
  assign n10287 = n10203 | n10286 ;
  assign n3710 = n3162 & n3701 ;
  assign n3077 = x[70] & n3031 ;
  assign n3103 = x[71] & n3096 ;
  assign n10182 = n3077 | n3103 ;
  assign n10183 = x[72] & n3027 ;
  assign n10184 = n10182 | n10183 ;
  assign n10185 = n3710 | n10184 ;
  assign n29712 = ~n10185 ;
  assign n10186 = x[41] & n29712 ;
  assign n10187 = n29184 & n10185 ;
  assign n10188 = n10186 | n10187 ;
  assign n9593 = n9589 & n9591 ;
  assign n9594 = n9556 | n9593 ;
  assign n9036 = n9027 & n9034 ;
  assign n6469 = n2321 & n6466 ;
  assign n2178 = n29619 & n2174 ;
  assign n29713 = ~n2177 ;
  assign n2179 = n29713 & n2178 ;
  assign n2215 = x[64] & n2179 ;
  assign n2260 = x[65] & n2244 ;
  assign n9037 = n2215 | n2260 ;
  assign n9038 = x[66] & n2175 ;
  assign n9039 = n9037 | n9038 ;
  assign n9040 = n6469 | n9039 ;
  assign n29714 = ~n9040 ;
  assign n9041 = x[47] & n29714 ;
  assign n9042 = n29621 & n9040 ;
  assign n9043 = n9041 | n9042 ;
  assign n29715 = ~n9043 ;
  assign n9044 = n9036 & n29715 ;
  assign n29716 = ~n9036 ;
  assign n9536 = n29716 & n9043 ;
  assign n9537 = n9044 | n9536 ;
  assign n6389 = n2635 & n6379 ;
  assign n2503 = x[67] & n2492 ;
  assign n2573 = x[68] & n2557 ;
  assign n9538 = n2503 | n2573 ;
  assign n9539 = x[69] & n2488 ;
  assign n9540 = n9538 | n9539 ;
  assign n9541 = n6389 | n9540 ;
  assign n29717 = ~n9541 ;
  assign n9542 = x[44] & n29717 ;
  assign n9543 = n29400 & n9541 ;
  assign n9544 = n9542 | n9543 ;
  assign n29718 = ~n9544 ;
  assign n9545 = n9537 & n29718 ;
  assign n29719 = ~n9537 ;
  assign n9595 = n29719 & n9544 ;
  assign n9596 = n9545 | n9595 ;
  assign n29720 = ~n9596 ;
  assign n9597 = n9594 & n29720 ;
  assign n29721 = ~n9594 ;
  assign n10189 = n29721 & n9596 ;
  assign n10190 = n9597 | n10189 ;
  assign n29722 = ~n10188 ;
  assign n10191 = n29722 & n10190 ;
  assign n29723 = ~n10190 ;
  assign n10288 = n10188 & n29723 ;
  assign n10289 = n10191 | n10288 ;
  assign n29724 = ~n10289 ;
  assign n10290 = n10287 & n29724 ;
  assign n29725 = ~n10287 ;
  assign n10904 = n29725 & n10289 ;
  assign n10905 = n10290 | n10904 ;
  assign n3576 = n3289 & n3574 ;
  assign n3457 = x[73] & n3443 ;
  assign n3547 = x[74] & n3508 ;
  assign n10906 = n3457 | n3547 ;
  assign n10907 = x[75] & n3439 ;
  assign n10908 = n10906 | n10907 ;
  assign n10909 = n3576 | n10908 ;
  assign n29726 = ~n10909 ;
  assign n10910 = x[38] & n29726 ;
  assign n10911 = n28996 & n10909 ;
  assign n10912 = n10910 | n10911 ;
  assign n10913 = n10905 | n10912 ;
  assign n10914 = n10905 & n10912 ;
  assign n29727 = ~n10914 ;
  assign n11054 = n10913 & n29727 ;
  assign n11055 = n11053 & n11054 ;
  assign n11472 = n11053 | n11054 ;
  assign n29728 = ~n11055 ;
  assign n11473 = n29728 & n11472 ;
  assign n29729 = ~n11471 ;
  assign n11662 = n29729 & n11473 ;
  assign n29730 = ~n11473 ;
  assign n12162 = n11471 & n29730 ;
  assign n12163 = n11662 | n12162 ;
  assign n12164 = n12161 | n12163 ;
  assign n12165 = n12161 & n12163 ;
  assign n29731 = ~n12165 ;
  assign n12259 = n12164 & n29731 ;
  assign n29732 = ~n12258 ;
  assign n12485 = n29732 & n12259 ;
  assign n29733 = ~n12259 ;
  assign n12486 = n12258 & n29733 ;
  assign n12487 = n12485 | n12486 ;
  assign n12884 = n12270 | n12883 ;
  assign n29734 = ~n12487 ;
  assign n12885 = n29734 & n12884 ;
  assign n29735 = ~n12884 ;
  assign n13114 = n12487 & n29735 ;
  assign n13115 = n12885 | n13114 ;
  assign n4644 = n1293 & n4632 ;
  assign n4538 = x[82] & n4514 ;
  assign n4596 = x[83] & n4572 ;
  assign n13116 = n4538 | n4596 ;
  assign n13117 = x[84] & n4504 ;
  assign n13118 = n13116 | n13117 ;
  assign n13119 = n4644 | n13118 ;
  assign n29736 = ~n13119 ;
  assign n13120 = x[29] & n29736 ;
  assign n13121 = n28483 & n13119 ;
  assign n13122 = n13120 | n13121 ;
  assign n29737 = ~n13122 ;
  assign n13125 = n13115 & n29737 ;
  assign n29738 = ~n13115 ;
  assign n13126 = n29738 & n13122 ;
  assign n13127 = n13125 | n13126 ;
  assign n13137 = n13128 & n13135 ;
  assign n13400 = n13152 & n13399 ;
  assign n13401 = n13153 | n13400 ;
  assign n13402 = n13142 & n13401 ;
  assign n13403 = n13137 | n13402 ;
  assign n13404 = n13127 | n13403 ;
  assign n13405 = n13127 & n13403 ;
  assign n29739 = ~n13405 ;
  assign n13850 = n13404 & n29739 ;
  assign n1523 = n452 & n1522 ;
  assign n348 = x[85] & n330 ;
  assign n395 = x[86] & n390 ;
  assign n13851 = n348 | n395 ;
  assign n13852 = x[87] & n322 ;
  assign n13853 = n13851 | n13852 ;
  assign n13854 = n1523 | n13853 ;
  assign n29740 = ~n13854 ;
  assign n13855 = x[26] & n29740 ;
  assign n13856 = n28342 & n13854 ;
  assign n13857 = n13855 | n13856 ;
  assign n13858 = n13850 & n13857 ;
  assign n13123 = n13115 | n13122 ;
  assign n13124 = n13115 & n13122 ;
  assign n29741 = ~n13124 ;
  assign n13759 = n13123 & n29741 ;
  assign n29742 = ~n13403 ;
  assign n13760 = n29742 & n13759 ;
  assign n29743 = ~n13759 ;
  assign n14684 = n13403 & n29743 ;
  assign n14685 = n13760 | n14684 ;
  assign n14686 = n13857 | n14685 ;
  assign n29744 = ~n13858 ;
  assign n14751 = n29744 & n14686 ;
  assign n29745 = ~n14751 ;
  assign n14752 = n14188 & n29745 ;
  assign n14687 = n13857 & n14685 ;
  assign n14688 = n13867 & n13870 ;
  assign n29746 = ~n13880 ;
  assign n13884 = n29746 & n13882 ;
  assign n29747 = ~n13882 ;
  assign n14691 = n13880 & n29747 ;
  assign n14692 = n13884 | n14691 ;
  assign n14745 = n14692 & n14743 ;
  assign n14746 = n13883 | n14745 ;
  assign n14747 = n14689 & n14746 ;
  assign n14748 = n14688 | n14747 ;
  assign n14749 = n14686 & n14748 ;
  assign n14750 = n14687 | n14749 ;
  assign n29748 = ~n14750 ;
  assign n14753 = n14686 & n29748 ;
  assign n14754 = n14752 | n14753 ;
  assign n5321 = n1482 & n5302 ;
  assign n5274 = x[88] & n5240 ;
  assign n6253 = x[89] & n6179 ;
  assign n14755 = n5274 | n6253 ;
  assign n14756 = x[90] & n5238 ;
  assign n14757 = n14755 | n14756 ;
  assign n14758 = n5321 | n14757 ;
  assign n29749 = ~n14758 ;
  assign n14759 = x[23] & n29749 ;
  assign n14760 = n28221 & n14758 ;
  assign n14761 = n14759 | n14760 ;
  assign n29750 = ~n14761 ;
  assign n14762 = n14754 & n29750 ;
  assign n29751 = ~n14754 ;
  assign n15526 = n29751 & n14761 ;
  assign n15527 = n14762 | n15526 ;
  assign n15528 = n15525 & n15527 ;
  assign n15697 = n15525 | n15527 ;
  assign n29752 = ~n15528 ;
  assign n15698 = n29752 & n15697 ;
  assign n15699 = n15696 & n15698 ;
  assign n16194 = n15696 | n15698 ;
  assign n29753 = ~n15699 ;
  assign n16195 = n29753 & n16194 ;
  assign n16196 = n16193 & n16195 ;
  assign n16698 = n16193 | n16195 ;
  assign n29754 = ~n16196 ;
  assign n16699 = n29754 & n16698 ;
  assign n16700 = n16697 & n16699 ;
  assign n17156 = n16697 | n16699 ;
  assign n29755 = ~n16700 ;
  assign n17483 = n29755 & n17156 ;
  assign n29756 = ~n17155 ;
  assign n17485 = n29756 & n17483 ;
  assign n29757 = ~n17483 ;
  assign n17659 = n17155 & n29757 ;
  assign n17660 = n17485 | n17659 ;
  assign n29758 = ~n17658 ;
  assign n17662 = n29758 & n17660 ;
  assign n29759 = ~n17660 ;
  assign n18697 = n17658 & n29759 ;
  assign n18698 = n17662 | n18697 ;
  assign n18748 = n17687 | n18747 ;
  assign n18749 = n18700 & n18748 ;
  assign n18750 = n17674 | n18749 ;
  assign n18751 = n18698 | n18750 ;
  assign n18753 = n18698 & n18750 ;
  assign n29760 = ~n18753 ;
  assign n18892 = n18751 & n29760 ;
  assign n12732 = n2867 & n12695 ;
  assign n12692 = x[100] & n12633 ;
  assign n14401 = x[101] & n13533 ;
  assign n18893 = n12692 | n14401 ;
  assign n18894 = x[102] & n12631 ;
  assign n18895 = n18893 | n18894 ;
  assign n18896 = n12732 | n18895 ;
  assign n29761 = ~n18896 ;
  assign n18897 = x[11] & n29761 ;
  assign n18898 = n27892 & n18896 ;
  assign n18899 = n18897 | n18898 ;
  assign n29762 = ~n18899 ;
  assign n18900 = n18892 & n29762 ;
  assign n29763 = ~n18892 ;
  assign n20050 = n29763 & n18899 ;
  assign n20051 = n18900 | n20050 ;
  assign n20052 = n18915 & n18918 ;
  assign n20089 = n18953 | n20088 ;
  assign n20090 = n20056 & n20089 ;
  assign n20091 = n18940 | n20090 ;
  assign n20092 = n19524 & n20091 ;
  assign n20093 = n19523 | n20092 ;
  assign n20094 = n20053 & n20093 ;
  assign n20095 = n20052 | n20094 ;
  assign n20096 = n20051 | n20095 ;
  assign n20098 = n20051 & n20095 ;
  assign n29764 = ~n20098 ;
  assign n20183 = n20096 & n29764 ;
  assign n15365 = n3409 & n15308 ;
  assign n15281 = x[103] & n15246 ;
  assign n17284 = x[104] & n16288 ;
  assign n20184 = n15281 | n17284 ;
  assign n20185 = x[105] & n15244 ;
  assign n20186 = n20184 | n20185 ;
  assign n20187 = n15365 | n20186 ;
  assign n29765 = ~n20187 ;
  assign n20188 = x[8] & n29765 ;
  assign n20189 = n27845 & n20187 ;
  assign n20190 = n20188 | n20189 ;
  assign n20872 = n20183 | n20190 ;
  assign n20191 = n20183 & n20190 ;
  assign n20873 = n20871 & n20872 ;
  assign n20874 = n20191 | n20873 ;
  assign n29766 = ~n20874 ;
  assign n20875 = n20872 & n29766 ;
  assign n17661 = n17658 & n17660 ;
  assign n17663 = n17658 | n17660 ;
  assign n29767 = ~n17661 ;
  assign n17664 = n29767 & n17663 ;
  assign n29768 = ~n18750 ;
  assign n18752 = n17664 & n29768 ;
  assign n29769 = ~n17664 ;
  assign n18902 = n29769 & n18750 ;
  assign n18903 = n18752 | n18902 ;
  assign n18904 = n18899 | n18903 ;
  assign n18905 = n18899 & n18903 ;
  assign n29770 = ~n18905 ;
  assign n18906 = n18904 & n29770 ;
  assign n29771 = ~n20095 ;
  assign n20097 = n18906 & n29771 ;
  assign n29772 = ~n18906 ;
  assign n21109 = n29772 & n20095 ;
  assign n21110 = n20097 | n21109 ;
  assign n21111 = n20190 & n21110 ;
  assign n29773 = ~n21111 ;
  assign n21112 = n20872 & n29773 ;
  assign n21281 = n20200 | n21113 ;
  assign n21282 = n21280 & n21281 ;
  assign n21283 = n21114 | n21282 ;
  assign n29774 = ~n21112 ;
  assign n21335 = n29774 & n21283 ;
  assign n21336 = n20875 | n21335 ;
  assign n18450 = n3876 & n18392 ;
  assign n18364 = x[106] & n18329 ;
  assign n18537 = x[107] & n18514 ;
  assign n21337 = n18364 | n18537 ;
  assign n21338 = x[108] & n18327 ;
  assign n21339 = n21337 | n21338 ;
  assign n21340 = n18450 | n21339 ;
  assign n29775 = ~n21340 ;
  assign n21341 = x[5] & n29775 ;
  assign n21342 = n27813 & n21340 ;
  assign n21343 = n21341 | n21342 ;
  assign n21344 = n21336 | n21343 ;
  assign n21345 = n21336 & n21343 ;
  assign n29776 = ~n21345 ;
  assign n22283 = n21344 & n29776 ;
  assign n22284 = n22282 & n22283 ;
  assign n22362 = n22282 | n22283 ;
  assign n29777 = ~n22284 ;
  assign n22363 = n29777 & n22362 ;
  assign n29778 = ~n22361 ;
  assign n22364 = n29778 & n22363 ;
  assign n29779 = ~n22363 ;
  assign n22366 = n22361 & n29779 ;
  assign n22367 = n22364 | n22366 ;
  assign n22377 = n22368 & n22375 ;
  assign n23037 = n22377 | n23036 ;
  assign n23038 = n22367 | n23037 ;
  assign n23039 = n22367 & n23037 ;
  assign n29780 = ~n23039 ;
  assign n176 = n23038 & n29780 ;
  assign n22365 = n22361 & n22363 ;
  assign n23040 = n22365 | n23039 ;
  assign n597 = n595 & n596 ;
  assign n598 = n27618 | n597 ;
  assign n24561 = x[111] & x[112] ;
  assign n599 = x[111] | x[112] ;
  assign n29781 = ~n24561 ;
  assign n4439 = n29781 & n599 ;
  assign n4440 = n598 & n4439 ;
  assign n4441 = n598 | n4439 ;
  assign n29782 = ~n4440 ;
  assign n4442 = n29782 & n4441 ;
  assign n19707 = n4442 & n19656 ;
  assign n19775 = x[110] & n19723 ;
  assign n19876 = x[111] & n19829 ;
  assign n22345 = n19775 | n19876 ;
  assign n22346 = x[112] & n19655 ;
  assign n22347 = n22345 | n22346 ;
  assign n22348 = n19707 | n22347 ;
  assign n22349 = x[2] | n22348 ;
  assign n22350 = x[2] & n22348 ;
  assign n29783 = ~n22350 ;
  assign n22351 = n22349 & n29783 ;
  assign n15368 = n3223 & n15308 ;
  assign n15298 = x[104] & n15246 ;
  assign n17329 = x[105] & n16288 ;
  assign n20174 = n15298 | n17329 ;
  assign n20175 = x[106] & n15244 ;
  assign n20176 = n20174 | n20175 ;
  assign n20177 = n15368 | n20176 ;
  assign n29784 = ~n20177 ;
  assign n20178 = x[8] & n29784 ;
  assign n20179 = n27845 & n20177 ;
  assign n20180 = n20178 | n20179 ;
  assign n18754 = n17661 | n18753 ;
  assign n17481 = n17152 & n17479 ;
  assign n17482 = n16710 | n17481 ;
  assign n17484 = n17482 & n17483 ;
  assign n17486 = n16700 | n17484 ;
  assign n8731 = n2438 & n8706 ;
  assign n8690 = x[95] & n8645 ;
  assign n9844 = x[96] & n9278 ;
  assign n16681 = n8690 | n9844 ;
  assign n16682 = x[97] & n8643 ;
  assign n16683 = n16681 | n16682 ;
  assign n16684 = n8731 | n16683 ;
  assign n29785 = ~n16684 ;
  assign n16685 = x[17] & n29785 ;
  assign n16686 = n28039 & n16684 ;
  assign n16687 = n16685 | n16686 ;
  assign n16197 = n15699 | n16196 ;
  assign n14763 = n14754 & n14761 ;
  assign n15529 = n14763 | n15528 ;
  assign n5337 = n2046 & n5302 ;
  assign n5255 = x[89] & n5240 ;
  assign n6237 = x[90] & n6179 ;
  assign n14674 = n5255 | n6237 ;
  assign n14675 = x[91] & n5238 ;
  assign n14676 = n14674 | n14675 ;
  assign n14677 = n5337 | n14676 ;
  assign n29786 = ~n14677 ;
  assign n14678 = x[23] & n29786 ;
  assign n14679 = n28221 & n14677 ;
  assign n14680 = n14678 | n14679 ;
  assign n14189 = n13850 | n13857 ;
  assign n14190 = n14188 & n14189 ;
  assign n14191 = n13858 | n14190 ;
  assign n4656 = n1239 & n4632 ;
  assign n4557 = x[83] & n4514 ;
  assign n4617 = x[84] & n4572 ;
  assign n13100 = n4557 | n4617 ;
  assign n13101 = x[85] & n4504 ;
  assign n13102 = n13100 | n13101 ;
  assign n13103 = n4656 | n13102 ;
  assign n29787 = ~n13103 ;
  assign n13104 = x[29] & n29787 ;
  assign n13105 = n28483 & n13103 ;
  assign n13106 = n13104 | n13105 ;
  assign n11474 = n11471 & n11473 ;
  assign n12166 = n11474 | n12165 ;
  assign n4049 = n1741 & n4041 ;
  assign n3927 = x[77] & n3910 ;
  assign n3982 = x[78] & n3975 ;
  assign n11453 = n3927 | n3982 ;
  assign n11454 = x[79] & n3906 ;
  assign n11455 = n11453 | n11454 ;
  assign n11456 = n4049 | n11455 ;
  assign n29788 = ~n11456 ;
  assign n11457 = x[35] & n29788 ;
  assign n11458 = n28822 & n11456 ;
  assign n11459 = n11457 | n11458 ;
  assign n11058 = n10914 | n11055 ;
  assign n3578 = n2750 & n3574 ;
  assign n3458 = x[74] & n3443 ;
  assign n3526 = x[75] & n3508 ;
  assign n10895 = n3458 | n3526 ;
  assign n10896 = x[76] & n3439 ;
  assign n10897 = n10895 | n10896 ;
  assign n10898 = n3578 | n10897 ;
  assign n29789 = ~n10898 ;
  assign n10899 = x[38] & n29789 ;
  assign n10900 = n28996 & n10898 ;
  assign n10901 = n10899 | n10900 ;
  assign n10192 = n10188 & n10190 ;
  assign n10291 = n10287 & n10289 ;
  assign n10292 = n10192 | n10291 ;
  assign n5982 = n2635 & n5976 ;
  assign n2537 = x[68] & n2492 ;
  assign n2576 = x[69] & n2557 ;
  assign n9524 = n2537 | n2576 ;
  assign n9525 = x[70] & n2488 ;
  assign n9526 = n9524 | n9525 ;
  assign n9527 = n5982 | n9526 ;
  assign n29790 = ~n9527 ;
  assign n9528 = x[44] & n29790 ;
  assign n9529 = n29400 & n9527 ;
  assign n9530 = n9528 | n9529 ;
  assign n27695 = x[47] & x[48] ;
  assign n1858 = x[47] | x[48] ;
  assign n29791 = ~n27695 ;
  assign n1859 = n29791 & n1858 ;
  assign n8396 = x[64] & n1859 ;
  assign n9045 = n9036 & n9043 ;
  assign n9046 = n8396 & n9045 ;
  assign n9047 = n8396 | n9045 ;
  assign n29792 = ~n9046 ;
  assign n9048 = n29792 & n9047 ;
  assign n6502 = n2321 & n6494 ;
  assign n2188 = x[65] & n2179 ;
  assign n2282 = x[66] & n2244 ;
  assign n9049 = n2188 | n2282 ;
  assign n9050 = x[67] & n2175 ;
  assign n9051 = n9049 | n9050 ;
  assign n9052 = n6502 | n9051 ;
  assign n29793 = ~n9052 ;
  assign n9053 = x[47] & n29793 ;
  assign n9054 = n29621 & n9052 ;
  assign n9055 = n9053 | n9054 ;
  assign n29794 = ~n9055 ;
  assign n9056 = n9048 & n29794 ;
  assign n29795 = ~n9048 ;
  assign n9531 = n29795 & n9055 ;
  assign n9532 = n9056 | n9531 ;
  assign n9533 = n9530 & n9532 ;
  assign n9534 = n9530 | n9532 ;
  assign n29796 = ~n9533 ;
  assign n9535 = n29796 & n9534 ;
  assign n9546 = n9537 & n9544 ;
  assign n9598 = n9594 & n9596 ;
  assign n9599 = n9546 | n9598 ;
  assign n29797 = ~n9599 ;
  assign n9600 = n9535 & n29797 ;
  assign n29798 = ~n9535 ;
  assign n10172 = n29798 & n9599 ;
  assign n10173 = n9600 | n10172 ;
  assign n3737 = n3162 & n3733 ;
  assign n3075 = x[71] & n3031 ;
  assign n3124 = x[72] & n3096 ;
  assign n10174 = n3075 | n3124 ;
  assign n10175 = x[73] & n3027 ;
  assign n10176 = n10174 | n10175 ;
  assign n10177 = n3737 | n10176 ;
  assign n29799 = ~n10177 ;
  assign n10178 = x[41] & n29799 ;
  assign n10179 = n29184 & n10177 ;
  assign n10180 = n10178 | n10179 ;
  assign n10181 = n10173 & n10180 ;
  assign n10293 = n10173 | n10180 ;
  assign n29800 = ~n10181 ;
  assign n10294 = n29800 & n10293 ;
  assign n29801 = ~n10292 ;
  assign n10878 = n29801 & n10294 ;
  assign n29802 = ~n10294 ;
  assign n10902 = n10292 & n29802 ;
  assign n10903 = n10878 | n10902 ;
  assign n29803 = ~n10903 ;
  assign n11056 = n10901 & n29803 ;
  assign n29804 = ~n10901 ;
  assign n11057 = n29804 & n10903 ;
  assign n11059 = n11056 | n11057 ;
  assign n11060 = n11058 & n11059 ;
  assign n11460 = n11057 | n11058 ;
  assign n11461 = n11056 | n11460 ;
  assign n29805 = ~n11060 ;
  assign n11462 = n29805 & n11461 ;
  assign n11463 = n11459 | n11462 ;
  assign n11464 = n11459 & n11462 ;
  assign n29806 = ~n11464 ;
  assign n12167 = n11463 & n29806 ;
  assign n12168 = n12166 & n12167 ;
  assign n12239 = n12166 | n12167 ;
  assign n29807 = ~n12168 ;
  assign n12240 = n29807 & n12239 ;
  assign n1005 = n779 & n1003 ;
  assign n710 = x[80] & n663 ;
  assign n761 = x[81] & n720 ;
  assign n12241 = n710 | n761 ;
  assign n12242 = x[82] & n652 ;
  assign n12243 = n12241 | n12242 ;
  assign n12244 = n1005 | n12243 ;
  assign n29808 = ~n12244 ;
  assign n12245 = x[32] & n29808 ;
  assign n12246 = n28658 & n12244 ;
  assign n12247 = n12245 | n12246 ;
  assign n12249 = n12240 & n12247 ;
  assign n12250 = n12240 | n12247 ;
  assign n29809 = ~n12249 ;
  assign n12251 = n29809 & n12250 ;
  assign n12260 = n12258 & n12259 ;
  assign n12886 = n12258 | n12259 ;
  assign n29810 = ~n12260 ;
  assign n12887 = n29810 & n12886 ;
  assign n12888 = n12884 & n12887 ;
  assign n12889 = n12260 | n12888 ;
  assign n29811 = ~n12889 ;
  assign n12891 = n12251 & n29811 ;
  assign n29812 = ~n12251 ;
  assign n13109 = n29812 & n12889 ;
  assign n13110 = n12891 | n13109 ;
  assign n13111 = n13106 | n13110 ;
  assign n13112 = n13106 & n13110 ;
  assign n29813 = ~n13112 ;
  assign n13113 = n13111 & n29813 ;
  assign n13801 = n13141 | n13800 ;
  assign n13802 = n13759 & n13801 ;
  assign n13803 = n13124 | n13802 ;
  assign n29814 = ~n13803 ;
  assign n13804 = n13113 & n29814 ;
  assign n29815 = ~n13113 ;
  assign n13839 = n29815 & n13803 ;
  assign n13840 = n13804 | n13839 ;
  assign n1721 = n452 & n1720 ;
  assign n337 = x[86] & n330 ;
  assign n435 = x[87] & n390 ;
  assign n13841 = n337 | n435 ;
  assign n13842 = x[88] & n322 ;
  assign n13843 = n13841 | n13842 ;
  assign n13844 = n1721 | n13843 ;
  assign n29816 = ~n13844 ;
  assign n13845 = x[26] & n29816 ;
  assign n13846 = n28342 & n13844 ;
  assign n13847 = n13845 | n13846 ;
  assign n13848 = n13840 | n13847 ;
  assign n13849 = n13840 & n13847 ;
  assign n29817 = ~n13849 ;
  assign n14192 = n13848 & n29817 ;
  assign n29818 = ~n14191 ;
  assign n14193 = n29818 & n14192 ;
  assign n29819 = ~n14192 ;
  assign n14681 = n14191 & n29819 ;
  assign n14682 = n14193 | n14681 ;
  assign n29820 = ~n14680 ;
  assign n15129 = n29820 & n14682 ;
  assign n29821 = ~n14682 ;
  assign n15530 = n14680 & n29821 ;
  assign n15531 = n15129 | n15530 ;
  assign n15532 = n15529 | n15531 ;
  assign n15533 = n15529 & n15531 ;
  assign n29822 = ~n15533 ;
  assign n15680 = n15532 & n29822 ;
  assign n7185 = n2410 & n7162 ;
  assign n7129 = x[92] & n7100 ;
  assign n7689 = x[93] & n7647 ;
  assign n15681 = n7129 | n7689 ;
  assign n15682 = x[94] & n7098 ;
  assign n15683 = n15681 | n15682 ;
  assign n15684 = n7185 | n15683 ;
  assign n29823 = ~n15684 ;
  assign n15685 = x[20] & n29823 ;
  assign n15686 = n28114 & n15684 ;
  assign n15687 = n15685 | n15686 ;
  assign n15688 = n15680 | n15687 ;
  assign n15689 = n15680 & n15687 ;
  assign n29824 = ~n15689 ;
  assign n16500 = n15688 & n29824 ;
  assign n29825 = ~n16197 ;
  assign n16502 = n29825 & n16500 ;
  assign n29826 = ~n16500 ;
  assign n16688 = n16197 & n29826 ;
  assign n16689 = n16502 | n16688 ;
  assign n29827 = ~n16687 ;
  assign n17159 = n29827 & n16689 ;
  assign n29828 = ~n16689 ;
  assign n17487 = n16687 & n29828 ;
  assign n17488 = n17159 | n17487 ;
  assign n17489 = n17486 | n17488 ;
  assign n17490 = n17486 & n17488 ;
  assign n29829 = ~n17490 ;
  assign n17642 = n17489 & n29829 ;
  assign n10584 = n2466 & n10542 ;
  assign n10500 = x[98] & n10481 ;
  assign n11874 = x[99] & n11232 ;
  assign n17643 = n10500 | n11874 ;
  assign n17644 = x[100] & n10479 ;
  assign n17645 = n17643 | n17644 ;
  assign n17646 = n10584 | n17645 ;
  assign n29830 = ~n17646 ;
  assign n17647 = x[14] & n29830 ;
  assign n17648 = n27956 & n17646 ;
  assign n17649 = n17647 | n17648 ;
  assign n17650 = n17642 | n17649 ;
  assign n17651 = n17642 & n17649 ;
  assign n29831 = ~n17651 ;
  assign n18755 = n17650 & n29831 ;
  assign n18756 = n18754 & n18755 ;
  assign n18878 = n18754 | n18755 ;
  assign n29832 = ~n18756 ;
  assign n18879 = n29832 & n18878 ;
  assign n12756 = n2626 & n12695 ;
  assign n12644 = x[101] & n12633 ;
  assign n14382 = x[102] & n13533 ;
  assign n18880 = n12644 | n14382 ;
  assign n18881 = x[103] & n12631 ;
  assign n18882 = n18880 | n18881 ;
  assign n18883 = n12756 | n18882 ;
  assign n29833 = ~n18883 ;
  assign n18884 = x[11] & n29833 ;
  assign n18885 = n27892 & n18883 ;
  assign n18886 = n18884 | n18885 ;
  assign n29834 = ~n18886 ;
  assign n18889 = n18879 & n29834 ;
  assign n29835 = ~n18879 ;
  assign n18890 = n29835 & n18886 ;
  assign n18891 = n18889 | n18890 ;
  assign n18901 = n18892 & n18899 ;
  assign n19530 = n18917 | n19529 ;
  assign n19531 = n18906 & n19530 ;
  assign n19532 = n18901 | n19531 ;
  assign n19533 = n18891 | n19532 ;
  assign n19534 = n18891 & n19532 ;
  assign n29836 = ~n19534 ;
  assign n20876 = n19533 & n29836 ;
  assign n29837 = ~n20180 ;
  assign n20877 = n29837 & n20876 ;
  assign n29838 = ~n20876 ;
  assign n20878 = n20180 & n29838 ;
  assign n20879 = n20877 | n20878 ;
  assign n21284 = n20190 | n21110 ;
  assign n21285 = n21283 & n21284 ;
  assign n21286 = n21111 | n21285 ;
  assign n29839 = ~n20879 ;
  assign n21287 = n29839 & n21286 ;
  assign n29840 = ~n21286 ;
  assign n21325 = n20879 & n29840 ;
  assign n21326 = n21287 | n21325 ;
  assign n18432 = n3639 & n18392 ;
  assign n18350 = x[107] & n18329 ;
  assign n18545 = x[108] & n18514 ;
  assign n21327 = n18350 | n18545 ;
  assign n21328 = x[109] & n18327 ;
  assign n21329 = n21327 | n21328 ;
  assign n21330 = n18432 | n21329 ;
  assign n29841 = ~n21330 ;
  assign n21331 = x[5] & n29841 ;
  assign n21332 = n27813 & n21330 ;
  assign n21333 = n21331 | n21332 ;
  assign n21334 = n21326 & n21333 ;
  assign n21998 = n21326 | n21333 ;
  assign n29842 = ~n21334 ;
  assign n21999 = n29842 & n21998 ;
  assign n22285 = n21345 | n22284 ;
  assign n29843 = ~n22285 ;
  assign n22286 = n21999 & n29843 ;
  assign n29844 = ~n21999 ;
  assign n22352 = n29844 & n22285 ;
  assign n22353 = n22286 | n22352 ;
  assign n22354 = n22351 & n22353 ;
  assign n23041 = n22351 | n22353 ;
  assign n29845 = ~n22354 ;
  assign n23042 = n29845 & n23041 ;
  assign n23043 = n23040 & n23042 ;
  assign n27693 = n23040 | n23042 ;
  assign n29846 = ~n23043 ;
  assign n177 = n29846 & n27693 ;
  assign n23044 = n22354 | n23043 ;
  assign n29847 = ~n21369 ;
  assign n21373 = n29847 & n21372 ;
  assign n29848 = ~n21372 ;
  assign n21374 = n21369 & n29848 ;
  assign n21375 = n21373 | n21374 ;
  assign n21992 = n21375 & n21991 ;
  assign n21993 = n21371 | n21992 ;
  assign n21994 = n21360 & n21993 ;
  assign n21995 = n21358 | n21994 ;
  assign n21996 = n21344 & n21995 ;
  assign n21997 = n21345 | n21996 ;
  assign n22000 = n21997 & n21999 ;
  assign n22001 = n21334 | n22000 ;
  assign n12716 = n3001 & n12695 ;
  assign n12688 = x[102] & n12633 ;
  assign n14376 = x[103] & n13533 ;
  assign n18864 = n12688 | n14376 ;
  assign n18865 = x[104] & n12631 ;
  assign n18866 = n18864 | n18865 ;
  assign n18867 = n12716 | n18866 ;
  assign n29849 = ~n18867 ;
  assign n18868 = x[11] & n29849 ;
  assign n18869 = n27892 & n18867 ;
  assign n18870 = n18868 | n18869 ;
  assign n10589 = n2977 & n10542 ;
  assign n10537 = x[99] & n10481 ;
  assign n11875 = x[100] & n11232 ;
  assign n17628 = n10537 | n11875 ;
  assign n17629 = x[101] & n10479 ;
  assign n17630 = n17628 | n17629 ;
  assign n17631 = n10589 | n17630 ;
  assign n29850 = ~n17631 ;
  assign n17632 = x[14] & n29850 ;
  assign n17633 = n27956 & n17631 ;
  assign n17634 = n17632 | n17633 ;
  assign n16690 = n16687 & n16689 ;
  assign n17157 = n17155 & n17156 ;
  assign n17158 = n16700 | n17157 ;
  assign n17160 = n16687 | n16689 ;
  assign n29851 = ~n16690 ;
  assign n17161 = n29851 & n17160 ;
  assign n17162 = n17158 & n17161 ;
  assign n17163 = n16690 | n17162 ;
  assign n5307 = n1841 & n5302 ;
  assign n5258 = x[90] & n5240 ;
  assign n6241 = x[91] & n6179 ;
  assign n14664 = n5258 | n6241 ;
  assign n14665 = x[92] & n5238 ;
  assign n14666 = n14664 | n14665 ;
  assign n14667 = n5307 | n14666 ;
  assign n29852 = ~n14667 ;
  assign n14668 = x[23] & n29852 ;
  assign n14669 = n28221 & n14667 ;
  assign n14670 = n14668 | n14669 ;
  assign n1454 = n452 & n1453 ;
  assign n339 = x[87] & n330 ;
  assign n431 = x[88] & n390 ;
  assign n13826 = n339 | n431 ;
  assign n13827 = x[89] & n322 ;
  assign n13828 = n13826 | n13827 ;
  assign n13829 = n1454 | n13828 ;
  assign n29853 = ~n13829 ;
  assign n13830 = x[26] & n29853 ;
  assign n13831 = n28342 & n13829 ;
  assign n13832 = n13830 | n13831 ;
  assign n4646 = n1213 & n4632 ;
  assign n4530 = x[84] & n4514 ;
  assign n4615 = x[85] & n4572 ;
  assign n13086 = n4530 | n4615 ;
  assign n13087 = x[86] & n4504 ;
  assign n13088 = n13086 | n13087 ;
  assign n13089 = n4646 | n13088 ;
  assign n29854 = ~n13089 ;
  assign n13090 = x[29] & n29854 ;
  assign n13091 = n28483 & n13089 ;
  assign n13092 = n13090 | n13091 ;
  assign n1058 = n779 & n1057 ;
  assign n696 = x[81] & n663 ;
  assign n749 = x[82] & n720 ;
  assign n12226 = n696 | n749 ;
  assign n12227 = x[83] & n652 ;
  assign n12228 = n12226 | n12227 ;
  assign n12229 = n1058 | n12228 ;
  assign n29855 = ~n12229 ;
  assign n12230 = x[32] & n29855 ;
  assign n12231 = n28658 & n12229 ;
  assign n12232 = n12230 | n12231 ;
  assign n4042 = n1270 & n4041 ;
  assign n3928 = x[78] & n3910 ;
  assign n3992 = x[79] & n3975 ;
  assign n11440 = n3928 | n3992 ;
  assign n11441 = x[80] & n3906 ;
  assign n11442 = n11440 | n11441 ;
  assign n11443 = n4042 | n11442 ;
  assign n29856 = ~n11443 ;
  assign n11444 = x[35] & n29856 ;
  assign n11445 = n28822 & n11443 ;
  assign n11446 = n11444 | n11445 ;
  assign n11061 = n10901 & n10903 ;
  assign n11062 = n11060 | n11061 ;
  assign n4800 = n2635 & n4790 ;
  assign n2496 = x[69] & n2492 ;
  assign n2578 = x[70] & n2557 ;
  assign n9511 = n2496 | n2578 ;
  assign n9512 = x[71] & n2488 ;
  assign n9513 = n9511 | n9512 ;
  assign n9514 = n4800 | n9513 ;
  assign n29857 = ~n9514 ;
  assign n9515 = x[44] & n29857 ;
  assign n9516 = n29400 & n9514 ;
  assign n9517 = n9515 | n9516 ;
  assign n9057 = n9048 & n9055 ;
  assign n9058 = n9046 | n9057 ;
  assign n6415 = n2321 & n6408 ;
  assign n2189 = x[66] & n2179 ;
  assign n2261 = x[67] & n2244 ;
  assign n9016 = n2189 | n2261 ;
  assign n9017 = x[68] & n2175 ;
  assign n9018 = n9016 | n9017 ;
  assign n9019 = n6415 | n9018 ;
  assign n9020 = x[47] | n9019 ;
  assign n9021 = x[47] & n9019 ;
  assign n29858 = ~n9021 ;
  assign n9022 = n9020 & n29858 ;
  assign n29859 = ~n8396 ;
  assign n8397 = x[50] & n29859 ;
  assign n27697 = x[49] & x[50] ;
  assign n1860 = x[49] | x[50] ;
  assign n29860 = ~n27697 ;
  assign n1861 = n29860 & n1860 ;
  assign n2007 = n1859 & n1861 ;
  assign n6443 = n2007 & n6437 ;
  assign n29861 = ~n1861 ;
  assign n1862 = n1859 & n29861 ;
  assign n8398 = x[65] & n1862 ;
  assign n27698 = x[48] & x[49] ;
  assign n1863 = x[48] | x[49] ;
  assign n29862 = ~n27698 ;
  assign n1864 = n29862 & n1863 ;
  assign n29863 = ~n1859 ;
  assign n1931 = n29863 & n1864 ;
  assign n8399 = x[64] & n1931 ;
  assign n8400 = n8398 | n8399 ;
  assign n8401 = n6443 | n8400 ;
  assign n29864 = ~n8401 ;
  assign n8402 = x[50] & n29864 ;
  assign n29865 = ~x[50] ;
  assign n8403 = n29865 & n8401 ;
  assign n8404 = n8402 | n8403 ;
  assign n29866 = ~n8404 ;
  assign n8405 = n8397 & n29866 ;
  assign n29867 = ~n8397 ;
  assign n9023 = n29867 & n8404 ;
  assign n9024 = n8405 | n9023 ;
  assign n9025 = n9022 & n9024 ;
  assign n9059 = n9022 | n9024 ;
  assign n29868 = ~n9025 ;
  assign n9060 = n29868 & n9059 ;
  assign n29869 = ~n9058 ;
  assign n9061 = n29869 & n9060 ;
  assign n29870 = ~n9060 ;
  assign n9518 = n9058 & n29870 ;
  assign n9519 = n9061 | n9518 ;
  assign n29871 = ~n9517 ;
  assign n9520 = n29871 & n9519 ;
  assign n29872 = ~n9519 ;
  assign n9522 = n9517 & n29872 ;
  assign n9523 = n9520 | n9522 ;
  assign n9601 = n9535 & n9599 ;
  assign n9602 = n9533 | n9601 ;
  assign n29873 = ~n9602 ;
  assign n9603 = n9523 & n29873 ;
  assign n29874 = ~n9523 ;
  assign n10162 = n29874 & n9602 ;
  assign n10163 = n9603 | n10162 ;
  assign n3176 = n2722 & n3162 ;
  assign n3048 = x[72] & n3031 ;
  assign n3149 = x[73] & n3096 ;
  assign n10164 = n3048 | n3149 ;
  assign n10165 = x[74] & n3027 ;
  assign n10166 = n10164 | n10165 ;
  assign n10167 = n3176 | n10166 ;
  assign n29875 = ~n10167 ;
  assign n10168 = x[41] & n29875 ;
  assign n10169 = n29184 & n10167 ;
  assign n10170 = n10168 | n10169 ;
  assign n10297 = n10163 | n10170 ;
  assign n10171 = n10163 & n10170 ;
  assign n10879 = n10292 & n10293 ;
  assign n10880 = n10181 | n10879 ;
  assign n10881 = n10297 & n10880 ;
  assign n10882 = n10171 | n10881 ;
  assign n29876 = ~n10882 ;
  assign n10883 = n10297 & n29876 ;
  assign n10295 = n10292 & n10294 ;
  assign n10296 = n10181 | n10295 ;
  assign n29877 = ~n10171 ;
  assign n10298 = n29877 & n10297 ;
  assign n29878 = ~n10298 ;
  assign n10884 = n10296 & n29878 ;
  assign n10885 = n10883 | n10884 ;
  assign n3600 = n1775 & n3574 ;
  assign n3464 = x[75] & n3443 ;
  assign n3523 = x[76] & n3508 ;
  assign n10886 = n3464 | n3523 ;
  assign n10887 = x[77] & n3439 ;
  assign n10888 = n10886 | n10887 ;
  assign n10889 = n3600 | n10888 ;
  assign n29879 = ~n10889 ;
  assign n10890 = x[38] & n29879 ;
  assign n10891 = n28996 & n10889 ;
  assign n10892 = n10890 | n10891 ;
  assign n10893 = n10885 | n10892 ;
  assign n10894 = n10885 & n10892 ;
  assign n29880 = ~n10894 ;
  assign n11063 = n10893 & n29880 ;
  assign n11064 = n11062 & n11063 ;
  assign n11447 = n11062 | n11063 ;
  assign n29881 = ~n11064 ;
  assign n11448 = n29881 & n11447 ;
  assign n29882 = ~n11446 ;
  assign n11450 = n29882 & n11448 ;
  assign n29883 = ~n11448 ;
  assign n12142 = n11446 & n29883 ;
  assign n12143 = n11450 | n12142 ;
  assign n12169 = n11464 | n12168 ;
  assign n12171 = n12143 | n12169 ;
  assign n12172 = n12143 & n12169 ;
  assign n29884 = ~n12172 ;
  assign n12235 = n12171 & n29884 ;
  assign n29885 = ~n12232 ;
  assign n12236 = n29885 & n12235 ;
  assign n29886 = ~n12235 ;
  assign n12237 = n12232 & n29886 ;
  assign n12238 = n12236 | n12237 ;
  assign n12466 = n12311 & n12465 ;
  assign n12468 = n12311 | n12465 ;
  assign n29887 = ~n12466 ;
  assign n12469 = n29887 & n12468 ;
  assign n12470 = n12463 & n12469 ;
  assign n12471 = n12314 | n12470 ;
  assign n12472 = n12303 & n12471 ;
  assign n12473 = n12304 | n12472 ;
  assign n12476 = n12473 & n12475 ;
  assign n12477 = n12293 | n12476 ;
  assign n12481 = n12477 & n12480 ;
  assign n12482 = n12283 | n12481 ;
  assign n12483 = n12273 & n12482 ;
  assign n12484 = n12270 | n12483 ;
  assign n12488 = n12484 & n12487 ;
  assign n12489 = n12260 | n12488 ;
  assign n12490 = n12251 & n12489 ;
  assign n12491 = n12249 | n12490 ;
  assign n12492 = n12238 | n12491 ;
  assign n12493 = n12238 & n12491 ;
  assign n29888 = ~n12493 ;
  assign n13095 = n12492 & n29888 ;
  assign n29889 = ~n13092 ;
  assign n13096 = n29889 & n13095 ;
  assign n29890 = ~n13095 ;
  assign n13097 = n13092 & n29890 ;
  assign n13098 = n13096 | n13097 ;
  assign n29891 = ~n12247 ;
  assign n12248 = n12240 & n29891 ;
  assign n29892 = ~n12240 ;
  assign n12861 = n29892 & n12247 ;
  assign n12862 = n12248 | n12861 ;
  assign n12890 = n12862 | n12889 ;
  assign n12892 = n12862 & n12889 ;
  assign n29893 = ~n12892 ;
  assign n13099 = n12890 & n29893 ;
  assign n13108 = n13099 & n13106 ;
  assign n13406 = n13124 | n13405 ;
  assign n13407 = n13113 & n13406 ;
  assign n13408 = n13108 | n13407 ;
  assign n13409 = n13098 | n13408 ;
  assign n13410 = n13098 & n13408 ;
  assign n29894 = ~n13410 ;
  assign n13835 = n13409 & n29894 ;
  assign n29895 = ~n13832 ;
  assign n13836 = n29895 & n13835 ;
  assign n29896 = ~n13835 ;
  assign n13837 = n13832 & n29896 ;
  assign n13838 = n13836 | n13837 ;
  assign n14194 = n14191 & n14192 ;
  assign n14195 = n13849 | n14194 ;
  assign n14196 = n13838 | n14195 ;
  assign n14197 = n13838 & n14195 ;
  assign n29897 = ~n14197 ;
  assign n15134 = n14196 & n29897 ;
  assign n29898 = ~n14670 ;
  assign n15135 = n29898 & n15134 ;
  assign n29899 = ~n15134 ;
  assign n15137 = n14670 & n29899 ;
  assign n15138 = n15135 | n15137 ;
  assign n14683 = n14680 & n14682 ;
  assign n15534 = n14683 | n15533 ;
  assign n29900 = ~n15138 ;
  assign n15535 = n29900 & n15534 ;
  assign n29901 = ~n15534 ;
  assign n15667 = n15138 & n29901 ;
  assign n15668 = n15535 | n15667 ;
  assign n7195 = n2152 & n7162 ;
  assign n7116 = x[93] & n7100 ;
  assign n7693 = x[94] & n7647 ;
  assign n15669 = n7116 | n7693 ;
  assign n15670 = x[95] & n7098 ;
  assign n15671 = n15669 | n15670 ;
  assign n15672 = n7195 | n15671 ;
  assign n29902 = ~n15672 ;
  assign n15673 = x[20] & n29902 ;
  assign n15674 = n28114 & n15672 ;
  assign n15675 = n15673 | n15674 ;
  assign n15677 = n15668 & n15675 ;
  assign n15678 = n15668 | n15675 ;
  assign n29903 = ~n15677 ;
  assign n15679 = n29903 & n15678 ;
  assign n16189 = n15706 & n16187 ;
  assign n16494 = n15706 | n16187 ;
  assign n29904 = ~n16189 ;
  assign n16495 = n29904 & n16494 ;
  assign n16496 = n16492 & n16495 ;
  assign n16497 = n15709 | n16496 ;
  assign n16498 = n16194 & n16497 ;
  assign n16499 = n15699 | n16498 ;
  assign n16501 = n16499 & n16500 ;
  assign n16503 = n15689 | n16501 ;
  assign n29905 = ~n16503 ;
  assign n16504 = n15679 & n29905 ;
  assign n29906 = ~n15679 ;
  assign n16666 = n29906 & n16503 ;
  assign n16667 = n16504 | n16666 ;
  assign n8732 = n2841 & n8706 ;
  assign n8680 = x[96] & n8645 ;
  assign n9873 = x[97] & n9278 ;
  assign n16668 = n8680 | n9873 ;
  assign n16669 = x[98] & n8643 ;
  assign n16670 = n16668 | n16669 ;
  assign n16671 = n8732 | n16670 ;
  assign n29907 = ~n16671 ;
  assign n16672 = x[17] & n29907 ;
  assign n16673 = n28039 & n16671 ;
  assign n16674 = n16672 | n16673 ;
  assign n16675 = n16667 | n16674 ;
  assign n16676 = n16667 & n16674 ;
  assign n29908 = ~n16676 ;
  assign n17452 = n16675 & n29908 ;
  assign n29909 = ~n17163 ;
  assign n17453 = n29909 & n17452 ;
  assign n29910 = ~n17452 ;
  assign n17637 = n17163 & n29910 ;
  assign n17638 = n17453 | n17637 ;
  assign n17639 = n17634 | n17638 ;
  assign n17640 = n17634 & n17638 ;
  assign n29911 = ~n17640 ;
  assign n17641 = n17639 & n29911 ;
  assign n18757 = n17651 | n18756 ;
  assign n29912 = ~n18757 ;
  assign n18759 = n17641 & n29912 ;
  assign n29913 = ~n17641 ;
  assign n18873 = n29913 & n18757 ;
  assign n18874 = n18759 | n18873 ;
  assign n18875 = n18870 | n18874 ;
  assign n18876 = n18870 & n18874 ;
  assign n29914 = ~n18876 ;
  assign n18877 = n18875 & n29914 ;
  assign n18888 = n18879 & n18886 ;
  assign n18887 = n18879 | n18886 ;
  assign n29915 = ~n18888 ;
  assign n20048 = n18887 & n29915 ;
  assign n20099 = n18905 | n20098 ;
  assign n20100 = n20048 & n20099 ;
  assign n20101 = n18888 | n20100 ;
  assign n29916 = ~n20101 ;
  assign n20102 = n18877 & n29916 ;
  assign n29917 = ~n18877 ;
  assign n20160 = n29917 & n20101 ;
  assign n20161 = n20102 | n20160 ;
  assign n15349 = n3199 & n15308 ;
  assign n15276 = x[105] & n15246 ;
  assign n17301 = x[106] & n16288 ;
  assign n20162 = n15276 | n17301 ;
  assign n20163 = x[107] & n15244 ;
  assign n20164 = n20162 | n20163 ;
  assign n20165 = n15349 | n20164 ;
  assign n29918 = ~n20165 ;
  assign n20166 = x[8] & n29918 ;
  assign n20167 = n27845 & n20165 ;
  assign n20168 = n20166 | n20167 ;
  assign n20169 = n20161 | n20168 ;
  assign n20170 = n20161 & n20168 ;
  assign n29919 = ~n20170 ;
  assign n20171 = n20169 & n29919 ;
  assign n21108 = n20180 & n20876 ;
  assign n29920 = ~n19532 ;
  assign n20049 = n29920 & n20048 ;
  assign n29921 = ~n20048 ;
  assign n20172 = n19532 & n29921 ;
  assign n20173 = n20049 | n20172 ;
  assign n20181 = n20173 | n20180 ;
  assign n20182 = n20173 & n20180 ;
  assign n29922 = ~n20182 ;
  assign n21288 = n20181 & n29922 ;
  assign n21289 = n21286 & n21288 ;
  assign n21290 = n21108 | n21289 ;
  assign n29923 = ~n21290 ;
  assign n21291 = n20171 & n29923 ;
  assign n29924 = ~n20171 ;
  assign n21309 = n29924 & n21290 ;
  assign n21310 = n21291 | n21309 ;
  assign n18447 = n3615 & n18392 ;
  assign n18374 = x[108] & n18329 ;
  assign n18533 = x[109] & n18514 ;
  assign n21311 = n18374 | n18533 ;
  assign n21312 = x[110] & n18327 ;
  assign n21313 = n21311 | n21312 ;
  assign n21314 = n18447 | n21313 ;
  assign n29925 = ~n21314 ;
  assign n21315 = x[5] & n29925 ;
  assign n21316 = n27813 & n21314 ;
  assign n21317 = n21315 | n21316 ;
  assign n21318 = n21310 | n21317 ;
  assign n21319 = n21310 & n21317 ;
  assign n29926 = ~n21319 ;
  assign n22097 = n21318 & n29926 ;
  assign n29927 = ~n22001 ;
  assign n22098 = n29927 & n22097 ;
  assign n29928 = ~n22097 ;
  assign n22334 = n22001 & n29928 ;
  assign n22335 = n22098 | n22334 ;
  assign n600 = n598 & n599 ;
  assign n601 = n24561 | n600 ;
  assign n27609 = x[112] & x[113] ;
  assign n602 = x[112] | x[113] ;
  assign n29929 = ~n27609 ;
  assign n4084 = n29929 & n602 ;
  assign n4085 = n601 | n4084 ;
  assign n4086 = n601 & n4084 ;
  assign n29930 = ~n4086 ;
  assign n4087 = n4085 & n29930 ;
  assign n19661 = n4087 & n19656 ;
  assign n19770 = x[111] & n19723 ;
  assign n19867 = x[112] & n19829 ;
  assign n22336 = n19770 | n19867 ;
  assign n22337 = x[113] & n19655 ;
  assign n22338 = n22336 | n22337 ;
  assign n22339 = n19661 | n22338 ;
  assign n29931 = ~n22339 ;
  assign n22340 = x[2] & n29931 ;
  assign n22341 = n27790 & n22339 ;
  assign n22342 = n22340 | n22341 ;
  assign n22343 = n22335 | n22342 ;
  assign n22344 = n22335 & n22342 ;
  assign n29932 = ~n22344 ;
  assign n23045 = n22343 & n29932 ;
  assign n23046 = n23044 | n23045 ;
  assign n23047 = n23044 & n23045 ;
  assign n29933 = ~n23047 ;
  assign n178 = n23046 & n29933 ;
  assign n21292 = n20171 & n21290 ;
  assign n21293 = n20170 | n21292 ;
  assign n29934 = ~n15675 ;
  assign n15676 = n15668 & n29934 ;
  assign n29935 = ~n15668 ;
  assign n16400 = n29935 & n15675 ;
  assign n16401 = n15676 | n16400 ;
  assign n16505 = n16401 | n16503 ;
  assign n16506 = n16401 & n16503 ;
  assign n29936 = ~n16506 ;
  assign n16677 = n16505 & n29936 ;
  assign n29937 = ~n16674 ;
  assign n16678 = n29937 & n16677 ;
  assign n29938 = ~n16677 ;
  assign n16679 = n16674 & n29938 ;
  assign n16680 = n16678 | n16679 ;
  assign n17164 = n16680 | n17163 ;
  assign n17165 = n16680 & n17163 ;
  assign n29939 = ~n17165 ;
  assign n17627 = n17164 & n29939 ;
  assign n29940 = ~n17634 ;
  assign n17635 = n17627 & n29940 ;
  assign n29941 = ~n17627 ;
  assign n18695 = n29941 & n17634 ;
  assign n18696 = n17635 | n18695 ;
  assign n18758 = n18696 | n18757 ;
  assign n18760 = n18696 & n18757 ;
  assign n29942 = ~n18760 ;
  assign n18863 = n18758 & n29942 ;
  assign n18872 = n18863 & n18870 ;
  assign n19535 = n18888 | n19534 ;
  assign n19536 = n18877 & n19535 ;
  assign n19537 = n18872 | n19536 ;
  assign n17636 = n17627 & n17634 ;
  assign n18233 = n17674 | n18232 ;
  assign n18234 = n17664 & n18233 ;
  assign n18235 = n17661 | n18234 ;
  assign n18236 = n17650 & n18235 ;
  assign n18237 = n17651 | n18236 ;
  assign n18238 = n17641 & n18237 ;
  assign n18239 = n17636 | n18238 ;
  assign n8766 = n2313 & n8706 ;
  assign n8681 = x[97] & n8645 ;
  assign n9846 = x[98] & n9278 ;
  assign n16653 = n8681 | n9846 ;
  assign n16654 = x[99] & n8643 ;
  assign n16655 = n16653 | n16654 ;
  assign n16656 = n8766 | n16655 ;
  assign n29943 = ~n16656 ;
  assign n16657 = x[17] & n29943 ;
  assign n16658 = n28039 & n16656 ;
  assign n16659 = n16657 | n16658 ;
  assign n16507 = n15677 | n16506 ;
  assign n7187 = n2000 & n7162 ;
  assign n7117 = x[94] & n7100 ;
  assign n7691 = x[95] & n7647 ;
  assign n15657 = n7117 | n7691 ;
  assign n15658 = x[96] & n7098 ;
  assign n15659 = n15657 | n15658 ;
  assign n15660 = n7187 | n15659 ;
  assign n29944 = ~n15660 ;
  assign n15661 = x[20] & n29944 ;
  assign n15662 = n28114 & n15660 ;
  assign n15663 = n15661 | n15662 ;
  assign n11449 = n11446 & n11448 ;
  assign n11451 = n11446 | n11448 ;
  assign n29945 = ~n11449 ;
  assign n11452 = n29945 & n11451 ;
  assign n29946 = ~n12169 ;
  assign n12170 = n11452 & n29946 ;
  assign n29947 = ~n11452 ;
  assign n12224 = n29947 & n12169 ;
  assign n12225 = n12170 | n12224 ;
  assign n12233 = n12225 | n12232 ;
  assign n12234 = n12225 & n12232 ;
  assign n29948 = ~n12234 ;
  assign n12859 = n12233 & n29948 ;
  assign n29949 = ~n12491 ;
  assign n12860 = n29949 & n12859 ;
  assign n29950 = ~n12859 ;
  assign n13084 = n12491 & n29950 ;
  assign n13085 = n12860 | n13084 ;
  assign n13093 = n13085 | n13092 ;
  assign n13094 = n13085 & n13092 ;
  assign n29951 = ~n13094 ;
  assign n13755 = n13093 & n29951 ;
  assign n29952 = ~n13408 ;
  assign n13756 = n29952 & n13755 ;
  assign n29953 = ~n13755 ;
  assign n13824 = n13408 & n29953 ;
  assign n13825 = n13756 | n13824 ;
  assign n13833 = n13825 | n13832 ;
  assign n13834 = n13825 & n13832 ;
  assign n29954 = ~n13834 ;
  assign n14591 = n13833 & n29954 ;
  assign n29955 = ~n14195 ;
  assign n14592 = n29955 & n14591 ;
  assign n29956 = ~n14591 ;
  assign n14671 = n14195 & n29956 ;
  assign n14672 = n14592 | n14671 ;
  assign n14673 = n14670 & n14672 ;
  assign n14773 = n14764 & n14771 ;
  assign n15124 = n14778 & n15123 ;
  assign n15125 = n14773 | n15124 ;
  assign n15126 = n14754 | n14761 ;
  assign n15127 = n15125 & n15126 ;
  assign n15128 = n14763 | n15127 ;
  assign n15130 = n14680 | n14682 ;
  assign n29957 = ~n14683 ;
  assign n15131 = n29957 & n15130 ;
  assign n15132 = n15128 & n15131 ;
  assign n15133 = n14683 | n15132 ;
  assign n15139 = n15133 & n15138 ;
  assign n15140 = n14673 | n15139 ;
  assign n5319 = n1685 & n5302 ;
  assign n5259 = x[91] & n5240 ;
  assign n6242 = x[92] & n6179 ;
  assign n14654 = n5259 | n6242 ;
  assign n14655 = x[93] & n5238 ;
  assign n14656 = n14654 | n14655 ;
  assign n14657 = n5319 | n14656 ;
  assign n29958 = ~n14657 ;
  assign n14658 = x[23] & n29958 ;
  assign n14659 = n28221 & n14657 ;
  assign n14660 = n14658 | n14659 ;
  assign n14198 = n13834 | n14197 ;
  assign n13411 = n13094 | n13410 ;
  assign n4051 = n1029 & n4041 ;
  assign n3931 = x[79] & n3910 ;
  assign n4015 = x[80] & n3975 ;
  assign n11431 = n3931 | n4015 ;
  assign n11432 = x[81] & n3906 ;
  assign n11433 = n11431 | n11432 ;
  assign n11434 = n4051 | n11433 ;
  assign n29959 = ~n11434 ;
  assign n11435 = x[35] & n29959 ;
  assign n11436 = n28822 & n11434 ;
  assign n11437 = n11435 | n11436 ;
  assign n11065 = n10894 | n11064 ;
  assign n3592 = n2084 & n3574 ;
  assign n3471 = x[76] & n3443 ;
  assign n3540 = x[77] & n3508 ;
  assign n10867 = n3471 | n3540 ;
  assign n10868 = x[78] & n3439 ;
  assign n10869 = n10867 | n10868 ;
  assign n10870 = n3592 | n10869 ;
  assign n29960 = ~n10870 ;
  assign n10871 = x[38] & n29960 ;
  assign n10872 = n28996 & n10870 ;
  assign n10873 = n10871 | n10872 ;
  assign n10299 = n10296 & n10297 ;
  assign n10300 = n10171 | n10299 ;
  assign n9521 = n9517 & n9519 ;
  assign n9604 = n9523 & n9602 ;
  assign n9605 = n9521 | n9604 ;
  assign n3706 = n2635 & n3701 ;
  assign n2519 = x[70] & n2492 ;
  assign n2585 = x[71] & n2557 ;
  assign n9500 = n2519 | n2585 ;
  assign n9501 = x[72] & n2488 ;
  assign n9502 = n9500 | n9501 ;
  assign n9503 = n3706 | n9502 ;
  assign n29961 = ~n9503 ;
  assign n9504 = x[44] & n29961 ;
  assign n9505 = n29400 & n9503 ;
  assign n9506 = n9504 | n9505 ;
  assign n9062 = n9058 & n9060 ;
  assign n9063 = n9025 | n9062 ;
  assign n8406 = n8397 & n8404 ;
  assign n6472 = n2007 & n6466 ;
  assign n1865 = n29863 & n1861 ;
  assign n29962 = ~n1864 ;
  assign n1866 = n29962 & n1865 ;
  assign n1891 = x[64] & n1866 ;
  assign n1949 = x[65] & n1931 ;
  assign n8407 = n1891 | n1949 ;
  assign n8408 = x[66] & n1862 ;
  assign n8409 = n8407 | n8408 ;
  assign n8410 = n6472 | n8409 ;
  assign n29963 = ~n8410 ;
  assign n8411 = x[50] & n29963 ;
  assign n8412 = n29865 & n8410 ;
  assign n8413 = n8411 | n8412 ;
  assign n29964 = ~n8413 ;
  assign n8414 = n8406 & n29964 ;
  assign n29965 = ~n8406 ;
  assign n9005 = n29965 & n8413 ;
  assign n9006 = n8414 | n9005 ;
  assign n6384 = n2321 & n6379 ;
  assign n2218 = x[67] & n2179 ;
  assign n2251 = x[68] & n2244 ;
  assign n9007 = n2218 | n2251 ;
  assign n9008 = x[69] & n2175 ;
  assign n9009 = n9007 | n9008 ;
  assign n9010 = n6384 | n9009 ;
  assign n29966 = ~n9010 ;
  assign n9011 = x[47] & n29966 ;
  assign n9012 = n29621 & n9010 ;
  assign n9013 = n9011 | n9012 ;
  assign n29967 = ~n9013 ;
  assign n9014 = n9006 & n29967 ;
  assign n29968 = ~n9006 ;
  assign n9064 = n29968 & n9013 ;
  assign n9065 = n9014 | n9064 ;
  assign n29969 = ~n9065 ;
  assign n9066 = n9063 & n29969 ;
  assign n29970 = ~n9063 ;
  assign n9507 = n29970 & n9065 ;
  assign n9508 = n9066 | n9507 ;
  assign n29971 = ~n9506 ;
  assign n9509 = n29971 & n9508 ;
  assign n29972 = ~n9508 ;
  assign n9606 = n9506 & n29972 ;
  assign n9607 = n9509 | n9606 ;
  assign n29973 = ~n9607 ;
  assign n9608 = n9605 & n29973 ;
  assign n29974 = ~n9605 ;
  assign n10151 = n29974 & n9607 ;
  assign n10152 = n9608 | n10151 ;
  assign n3291 = n3162 & n3289 ;
  assign n3059 = x[73] & n3031 ;
  assign n3145 = x[74] & n3096 ;
  assign n10153 = n3059 | n3145 ;
  assign n10154 = x[75] & n3027 ;
  assign n10155 = n10153 | n10154 ;
  assign n10156 = n3291 | n10155 ;
  assign n29975 = ~n10156 ;
  assign n10157 = x[41] & n29975 ;
  assign n10158 = n29184 & n10156 ;
  assign n10159 = n10157 | n10158 ;
  assign n10160 = n10152 | n10159 ;
  assign n10161 = n10152 & n10159 ;
  assign n29976 = ~n10161 ;
  assign n10301 = n10160 & n29976 ;
  assign n10302 = n10300 & n10301 ;
  assign n10874 = n10300 | n10301 ;
  assign n29977 = ~n10302 ;
  assign n10875 = n29977 & n10874 ;
  assign n29978 = ~n10873 ;
  assign n10876 = n29978 & n10875 ;
  assign n29979 = ~n10875 ;
  assign n11066 = n10873 & n29979 ;
  assign n11067 = n10876 | n11066 ;
  assign n11068 = n11065 | n11067 ;
  assign n11069 = n11065 & n11067 ;
  assign n29980 = ~n11069 ;
  assign n11438 = n11068 & n29980 ;
  assign n29981 = ~n11437 ;
  assign n11671 = n29981 & n11438 ;
  assign n29982 = ~n11438 ;
  assign n11672 = n11437 & n29982 ;
  assign n11673 = n11671 | n11672 ;
  assign n12173 = n11449 | n12172 ;
  assign n29983 = ~n11673 ;
  assign n12174 = n29983 & n12173 ;
  assign n29984 = ~n12173 ;
  assign n12211 = n11673 & n29984 ;
  assign n12212 = n12174 | n12211 ;
  assign n1295 = n779 & n1293 ;
  assign n709 = x[82] & n663 ;
  assign n760 = x[83] & n720 ;
  assign n12213 = n709 | n760 ;
  assign n12214 = x[84] & n652 ;
  assign n12215 = n12213 | n12214 ;
  assign n12216 = n1295 | n12215 ;
  assign n29985 = ~n12216 ;
  assign n12217 = x[32] & n29985 ;
  assign n12218 = n28658 & n12216 ;
  assign n12219 = n12217 | n12218 ;
  assign n29986 = ~n12219 ;
  assign n12220 = n12212 & n29986 ;
  assign n29987 = ~n12212 ;
  assign n12856 = n29987 & n12219 ;
  assign n12857 = n12220 | n12856 ;
  assign n12858 = n12232 & n12235 ;
  assign n12893 = n12249 | n12892 ;
  assign n12894 = n12859 & n12893 ;
  assign n12895 = n12858 | n12894 ;
  assign n12896 = n12857 | n12895 ;
  assign n12898 = n12857 & n12895 ;
  assign n29988 = ~n12898 ;
  assign n13075 = n12896 & n29988 ;
  assign n4647 = n1522 & n4632 ;
  assign n4555 = x[85] & n4514 ;
  assign n4613 = x[86] & n4572 ;
  assign n13076 = n4555 | n4613 ;
  assign n13077 = x[87] & n4504 ;
  assign n13078 = n13076 | n13077 ;
  assign n13079 = n4647 | n13078 ;
  assign n29989 = ~n13079 ;
  assign n13080 = x[29] & n29989 ;
  assign n13081 = n28483 & n13079 ;
  assign n13082 = n13080 | n13081 ;
  assign n13083 = n13075 & n13082 ;
  assign n12221 = n12212 & n12219 ;
  assign n12222 = n12212 | n12219 ;
  assign n29990 = ~n12221 ;
  assign n12223 = n29990 & n12222 ;
  assign n29991 = ~n12895 ;
  assign n12897 = n12223 & n29991 ;
  assign n29992 = ~n12223 ;
  assign n13750 = n29992 & n12895 ;
  assign n13751 = n12897 | n13750 ;
  assign n13752 = n13082 | n13751 ;
  assign n29993 = ~n13083 ;
  assign n13811 = n29993 & n13752 ;
  assign n29994 = ~n13811 ;
  assign n13812 = n13411 & n29994 ;
  assign n13753 = n13082 & n13751 ;
  assign n13754 = n13092 & n13095 ;
  assign n29995 = ~n13106 ;
  assign n13107 = n13099 & n29995 ;
  assign n29996 = ~n13099 ;
  assign n13757 = n29996 & n13106 ;
  assign n13758 = n13107 | n13757 ;
  assign n13805 = n13758 & n13803 ;
  assign n13806 = n13112 | n13805 ;
  assign n13807 = n13755 & n13806 ;
  assign n13808 = n13754 | n13807 ;
  assign n13809 = n13752 & n13808 ;
  assign n13810 = n13753 | n13809 ;
  assign n29997 = ~n13810 ;
  assign n13813 = n13752 & n29997 ;
  assign n13814 = n13812 | n13813 ;
  assign n1485 = n452 & n1482 ;
  assign n334 = x[88] & n330 ;
  assign n405 = x[89] & n390 ;
  assign n13815 = n334 | n405 ;
  assign n13816 = x[90] & n322 ;
  assign n13817 = n13815 | n13816 ;
  assign n13818 = n1485 | n13817 ;
  assign n29998 = ~n13818 ;
  assign n13819 = x[26] & n29998 ;
  assign n13820 = n28342 & n13818 ;
  assign n13821 = n13819 | n13820 ;
  assign n29999 = ~n13821 ;
  assign n13822 = n13814 & n29999 ;
  assign n30000 = ~n13814 ;
  assign n14199 = n30000 & n13821 ;
  assign n14200 = n13822 | n14199 ;
  assign n14201 = n14198 & n14200 ;
  assign n14661 = n14198 | n14200 ;
  assign n30001 = ~n14201 ;
  assign n14662 = n30001 & n14661 ;
  assign n14663 = n14660 & n14662 ;
  assign n15141 = n14660 | n14662 ;
  assign n30002 = ~n14663 ;
  assign n15142 = n30002 & n15141 ;
  assign n15143 = n15140 & n15142 ;
  assign n15664 = n15140 | n15142 ;
  assign n30003 = ~n15143 ;
  assign n15665 = n30003 & n15664 ;
  assign n15666 = n15663 & n15665 ;
  assign n16202 = n15663 | n15665 ;
  assign n30004 = ~n15666 ;
  assign n16508 = n30004 & n16202 ;
  assign n16509 = n16507 & n16508 ;
  assign n16660 = n16507 | n16508 ;
  assign n30005 = ~n16509 ;
  assign n16661 = n30005 & n16660 ;
  assign n16662 = n16659 & n16661 ;
  assign n16664 = n16659 | n16661 ;
  assign n30006 = ~n16662 ;
  assign n16665 = n30006 & n16664 ;
  assign n17451 = n16674 & n16677 ;
  assign n17491 = n16690 | n17490 ;
  assign n17492 = n17452 & n17491 ;
  assign n17493 = n17451 | n17492 ;
  assign n30007 = ~n17493 ;
  assign n17494 = n16665 & n30007 ;
  assign n30008 = ~n16665 ;
  assign n17612 = n30008 & n17493 ;
  assign n17613 = n17494 | n17612 ;
  assign n10591 = n2867 & n10542 ;
  assign n10534 = x[100] & n10481 ;
  assign n11886 = x[101] & n11232 ;
  assign n17614 = n10534 | n11886 ;
  assign n17615 = x[102] & n10479 ;
  assign n17616 = n17614 | n17615 ;
  assign n17617 = n10591 | n17616 ;
  assign n30009 = ~n17617 ;
  assign n17618 = x[14] & n30009 ;
  assign n17619 = n27956 & n17617 ;
  assign n17620 = n17618 | n17619 ;
  assign n17621 = n17613 | n17620 ;
  assign n17622 = n17613 & n17620 ;
  assign n30010 = ~n17622 ;
  assign n18693 = n17621 & n30010 ;
  assign n30011 = ~n18239 ;
  assign n18694 = n30011 & n18693 ;
  assign n30012 = ~n18693 ;
  assign n18848 = n18239 & n30012 ;
  assign n18849 = n18694 | n18848 ;
  assign n12745 = n3409 & n12695 ;
  assign n12661 = x[103] & n12633 ;
  assign n14400 = x[104] & n13533 ;
  assign n18850 = n12661 | n14400 ;
  assign n18851 = x[105] & n12631 ;
  assign n18852 = n18850 | n18851 ;
  assign n18853 = n12745 | n18852 ;
  assign n30013 = ~n18853 ;
  assign n18854 = x[11] & n30013 ;
  assign n18855 = n27892 & n18853 ;
  assign n18856 = n18854 | n18855 ;
  assign n18857 = n18849 | n18856 ;
  assign n18858 = n18849 & n18856 ;
  assign n30014 = ~n18858 ;
  assign n20044 = n18857 & n30014 ;
  assign n30015 = ~n19537 ;
  assign n20045 = n30015 & n20044 ;
  assign n30016 = ~n20044 ;
  assign n20150 = n19537 & n30016 ;
  assign n20151 = n20045 | n20150 ;
  assign n15314 = n3876 & n15308 ;
  assign n15297 = x[106] & n15246 ;
  assign n17328 = x[107] & n16288 ;
  assign n20152 = n15297 | n17328 ;
  assign n20153 = x[108] & n15244 ;
  assign n20154 = n20152 | n20153 ;
  assign n20155 = n15314 | n20154 ;
  assign n30017 = ~n20155 ;
  assign n20156 = x[8] & n30017 ;
  assign n20157 = n27845 & n20155 ;
  assign n20158 = n20156 | n20157 ;
  assign n20159 = n20151 & n20158 ;
  assign n20884 = n20151 | n20158 ;
  assign n30018 = ~n20159 ;
  assign n21294 = n30018 & n20884 ;
  assign n30019 = ~n21294 ;
  assign n21295 = n21293 & n30019 ;
  assign n20880 = n20874 & n20879 ;
  assign n20881 = n20182 | n20880 ;
  assign n20882 = n20171 & n20881 ;
  assign n20883 = n20170 | n20882 ;
  assign n20885 = n20883 & n20884 ;
  assign n20886 = n20159 | n20885 ;
  assign n30020 = ~n20886 ;
  assign n21296 = n20884 & n30020 ;
  assign n21297 = n21295 | n21296 ;
  assign n18426 = n4246 & n18392 ;
  assign n18377 = x[109] & n18329 ;
  assign n18566 = x[110] & n18514 ;
  assign n21298 = n18377 | n18566 ;
  assign n21299 = x[111] & n18327 ;
  assign n21300 = n21298 | n21299 ;
  assign n21301 = n18426 | n21300 ;
  assign n30021 = ~n21301 ;
  assign n21302 = x[5] & n30021 ;
  assign n21303 = n27813 & n21301 ;
  assign n21304 = n21302 | n21303 ;
  assign n30022 = ~n21304 ;
  assign n21305 = n21297 & n30022 ;
  assign n30023 = ~n21297 ;
  assign n21307 = n30023 & n21304 ;
  assign n21308 = n21305 | n21307 ;
  assign n21320 = n20171 | n20881 ;
  assign n30024 = ~n20882 ;
  assign n21321 = n30024 & n21320 ;
  assign n22096 = n21317 & n21321 ;
  assign n22287 = n21998 & n22285 ;
  assign n22288 = n21334 | n22287 ;
  assign n22289 = n22097 & n22288 ;
  assign n22290 = n22096 | n22289 ;
  assign n22291 = n21308 | n22290 ;
  assign n22292 = n21308 & n22290 ;
  assign n30025 = ~n22292 ;
  assign n22322 = n22291 & n30025 ;
  assign n603 = n601 & n602 ;
  assign n604 = n27609 | n603 ;
  assign n24381 = x[113] & x[114] ;
  assign n605 = x[113] | x[114] ;
  assign n30026 = ~n24381 ;
  assign n4273 = n30026 & n605 ;
  assign n4274 = n604 & n4273 ;
  assign n4275 = n604 | n4273 ;
  assign n30027 = ~n4274 ;
  assign n4276 = n30027 & n4275 ;
  assign n19706 = n4276 & n19656 ;
  assign n19726 = x[112] & n19723 ;
  assign n19878 = x[113] & n19829 ;
  assign n22323 = n19726 | n19878 ;
  assign n22324 = x[114] & n19655 ;
  assign n22325 = n22323 | n22324 ;
  assign n22326 = n19706 | n22325 ;
  assign n30028 = ~n22326 ;
  assign n22327 = x[2] & n30028 ;
  assign n22328 = n27790 & n22326 ;
  assign n22329 = n22327 | n22328 ;
  assign n30029 = ~n22329 ;
  assign n22330 = n22322 & n30029 ;
  assign n30030 = ~n22322 ;
  assign n22332 = n30030 & n22329 ;
  assign n22333 = n22330 | n22332 ;
  assign n23048 = n22344 | n23047 ;
  assign n23049 = n22333 & n23048 ;
  assign n27696 = n22333 | n23048 ;
  assign n30031 = ~n23049 ;
  assign n179 = n30031 & n27696 ;
  assign n22331 = n22322 & n22329 ;
  assign n23050 = n22331 | n23049 ;
  assign n606 = n604 & n605 ;
  assign n607 = n24381 | n606 ;
  assign n27592 = x[114] & x[115] ;
  assign n608 = x[114] | x[115] ;
  assign n30032 = ~n27592 ;
  assign n4471 = n30032 & n608 ;
  assign n4472 = n607 | n4471 ;
  assign n4473 = n607 & n4471 ;
  assign n30033 = ~n4473 ;
  assign n4474 = n4472 & n30033 ;
  assign n19686 = n4474 & n19656 ;
  assign n19776 = x[113] & n19723 ;
  assign n19857 = x[114] & n19829 ;
  assign n22311 = n19776 | n19857 ;
  assign n22312 = x[115] & n19655 ;
  assign n22313 = n22311 | n22312 ;
  assign n22314 = n19686 | n22313 ;
  assign n30034 = ~n22314 ;
  assign n22315 = x[2] & n30034 ;
  assign n22316 = n27790 & n22314 ;
  assign n22317 = n22315 | n22316 ;
  assign n21306 = n21297 & n21304 ;
  assign n22293 = n21306 | n22292 ;
  assign n15364 = n3639 & n15308 ;
  assign n15253 = x[107] & n15246 ;
  assign n17326 = x[108] & n16288 ;
  assign n20140 = n15253 | n17326 ;
  assign n20141 = x[109] & n15244 ;
  assign n20142 = n20140 | n20141 ;
  assign n20143 = n15364 | n20142 ;
  assign n30035 = ~n20143 ;
  assign n20144 = x[8] & n30035 ;
  assign n20145 = n27845 & n20143 ;
  assign n20146 = n20144 | n20145 ;
  assign n30036 = ~n16659 ;
  assign n16663 = n30036 & n16661 ;
  assign n30037 = ~n16661 ;
  assign n17449 = n16659 & n30037 ;
  assign n17450 = n16663 | n17449 ;
  assign n17496 = n17450 & n17493 ;
  assign n17497 = n16662 | n17496 ;
  assign n16510 = n15666 | n16509 ;
  assign n7208 = n2438 & n7162 ;
  assign n7118 = x[95] & n7100 ;
  assign n7729 = x[96] & n7647 ;
  assign n15647 = n7118 | n7729 ;
  assign n15648 = x[97] & n7098 ;
  assign n15649 = n15647 | n15648 ;
  assign n15650 = n7208 | n15649 ;
  assign n30038 = ~n15650 ;
  assign n15651 = x[20] & n30038 ;
  assign n15652 = n28114 & n15650 ;
  assign n15653 = n15651 | n15652 ;
  assign n15144 = n14663 | n15143 ;
  assign n13823 = n13814 & n13821 ;
  assign n14202 = n13823 | n14201 ;
  assign n2048 = n452 & n2046 ;
  assign n349 = x[89] & n330 ;
  assign n434 = x[90] & n390 ;
  assign n13740 = n349 | n434 ;
  assign n13741 = x[91] & n322 ;
  assign n13742 = n13740 | n13741 ;
  assign n13743 = n2048 | n13742 ;
  assign n30039 = ~n13743 ;
  assign n13744 = x[26] & n30039 ;
  assign n13745 = n28342 & n13743 ;
  assign n13746 = n13744 | n13745 ;
  assign n13412 = n13075 | n13082 ;
  assign n13413 = n13411 & n13412 ;
  assign n13414 = n13083 | n13413 ;
  assign n12494 = n12234 | n12493 ;
  assign n12495 = n12223 & n12494 ;
  assign n12496 = n12221 | n12495 ;
  assign n4052 = n1003 & n4041 ;
  assign n3959 = x[80] & n3910 ;
  assign n3994 = x[81] & n3975 ;
  assign n11421 = n3959 | n3994 ;
  assign n11422 = x[82] & n3906 ;
  assign n11423 = n11421 | n11422 ;
  assign n11424 = n4052 | n11423 ;
  assign n30040 = ~n11424 ;
  assign n11425 = x[35] & n30040 ;
  assign n11426 = n28822 & n11424 ;
  assign n11427 = n11425 | n11426 ;
  assign n10877 = n10873 & n10875 ;
  assign n11070 = n10877 | n11069 ;
  assign n3580 = n1741 & n3574 ;
  assign n3476 = x[77] & n3443 ;
  assign n3545 = x[78] & n3508 ;
  assign n10855 = n3476 | n3545 ;
  assign n10856 = x[79] & n3439 ;
  assign n10857 = n10855 | n10856 ;
  assign n10858 = n3580 | n10857 ;
  assign n30041 = ~n10858 ;
  assign n10859 = x[38] & n30041 ;
  assign n10860 = n28996 & n10858 ;
  assign n10861 = n10859 | n10860 ;
  assign n10303 = n10161 | n10302 ;
  assign n3167 = n2750 & n3162 ;
  assign n3049 = x[74] & n3031 ;
  assign n3116 = x[75] & n3096 ;
  assign n10141 = n3049 | n3116 ;
  assign n10142 = x[76] & n3027 ;
  assign n10143 = n10141 | n10142 ;
  assign n10144 = n3167 | n10143 ;
  assign n30042 = ~n10144 ;
  assign n10145 = x[41] & n30042 ;
  assign n10146 = n29184 & n10144 ;
  assign n10147 = n10145 | n10146 ;
  assign n9510 = n9506 & n9508 ;
  assign n9609 = n9605 & n9607 ;
  assign n9610 = n9510 | n9609 ;
  assign n5989 = n2321 & n5976 ;
  assign n2191 = x[68] & n2179 ;
  assign n2271 = x[69] & n2244 ;
  assign n8993 = n2191 | n2271 ;
  assign n8994 = x[70] & n2175 ;
  assign n8995 = n8993 | n8994 ;
  assign n8996 = n5989 | n8995 ;
  assign n30043 = ~n8996 ;
  assign n8997 = x[47] & n30043 ;
  assign n8998 = n29621 & n8996 ;
  assign n8999 = n8997 | n8998 ;
  assign n27686 = x[50] & x[51] ;
  assign n1543 = x[50] | x[51] ;
  assign n30044 = ~n27686 ;
  assign n1544 = n30044 & n1543 ;
  assign n7914 = x[64] & n1544 ;
  assign n8415 = n8406 & n8413 ;
  assign n8416 = n7914 & n8415 ;
  assign n8417 = n7914 | n8415 ;
  assign n30045 = ~n8416 ;
  assign n8418 = n30045 & n8417 ;
  assign n6503 = n2007 & n6494 ;
  assign n1879 = x[65] & n1866 ;
  assign n1965 = x[66] & n1931 ;
  assign n8419 = n1879 | n1965 ;
  assign n8420 = x[67] & n1862 ;
  assign n8421 = n8419 | n8420 ;
  assign n8422 = n6503 | n8421 ;
  assign n30046 = ~n8422 ;
  assign n8423 = x[50] & n30046 ;
  assign n8424 = n29865 & n8422 ;
  assign n8425 = n8423 | n8424 ;
  assign n30047 = ~n8425 ;
  assign n8426 = n8418 & n30047 ;
  assign n30048 = ~n8418 ;
  assign n9000 = n30048 & n8425 ;
  assign n9001 = n8426 | n9000 ;
  assign n9002 = n8999 & n9001 ;
  assign n9003 = n8999 | n9001 ;
  assign n30049 = ~n9002 ;
  assign n9004 = n30049 & n9003 ;
  assign n9015 = n9006 & n9013 ;
  assign n9067 = n9063 & n9065 ;
  assign n9068 = n9015 | n9067 ;
  assign n30050 = ~n9068 ;
  assign n9069 = n9004 & n30050 ;
  assign n30051 = ~n9004 ;
  assign n9489 = n30051 & n9068 ;
  assign n9490 = n9069 | n9489 ;
  assign n3741 = n2635 & n3733 ;
  assign n2504 = x[71] & n2492 ;
  assign n2580 = x[72] & n2557 ;
  assign n9491 = n2504 | n2580 ;
  assign n9492 = x[73] & n2488 ;
  assign n9493 = n9491 | n9492 ;
  assign n9494 = n3741 | n9493 ;
  assign n30052 = ~n9494 ;
  assign n9495 = x[44] & n30052 ;
  assign n9496 = n29400 & n9494 ;
  assign n9497 = n9495 | n9496 ;
  assign n9498 = n9490 | n9497 ;
  assign n9499 = n9490 & n9497 ;
  assign n30053 = ~n9499 ;
  assign n9611 = n9498 & n30053 ;
  assign n30054 = ~n9610 ;
  assign n9612 = n30054 & n9611 ;
  assign n30055 = ~n9611 ;
  assign n10148 = n9610 & n30055 ;
  assign n10149 = n9612 | n10148 ;
  assign n30056 = ~n10149 ;
  assign n10304 = n10147 & n30056 ;
  assign n30057 = ~n10147 ;
  assign n10305 = n30057 & n10149 ;
  assign n10306 = n10304 | n10305 ;
  assign n10307 = n10303 & n10306 ;
  assign n10862 = n10303 | n10305 ;
  assign n10863 = n10304 | n10862 ;
  assign n30058 = ~n10307 ;
  assign n10864 = n30058 & n10863 ;
  assign n10865 = n10861 | n10864 ;
  assign n10866 = n10861 & n10864 ;
  assign n30059 = ~n10866 ;
  assign n11071 = n10865 & n30059 ;
  assign n11072 = n11070 & n11071 ;
  assign n11428 = n11070 | n11071 ;
  assign n30060 = ~n11072 ;
  assign n11429 = n30060 & n11428 ;
  assign n11430 = n11427 & n11429 ;
  assign n11676 = n11427 | n11429 ;
  assign n30061 = ~n11430 ;
  assign n11677 = n30061 & n11676 ;
  assign n11439 = n11437 & n11438 ;
  assign n12175 = n11437 | n11438 ;
  assign n30062 = ~n11439 ;
  assign n12176 = n30062 & n12175 ;
  assign n12177 = n12173 & n12176 ;
  assign n12178 = n11439 | n12177 ;
  assign n30063 = ~n12178 ;
  assign n12179 = n11677 & n30063 ;
  assign n30064 = ~n11677 ;
  assign n12197 = n30064 & n12178 ;
  assign n12198 = n12179 | n12197 ;
  assign n1240 = n779 & n1239 ;
  assign n708 = x[83] & n663 ;
  assign n759 = x[84] & n720 ;
  assign n12199 = n708 | n759 ;
  assign n12200 = x[85] & n652 ;
  assign n12201 = n12199 | n12200 ;
  assign n12202 = n1240 | n12201 ;
  assign n30065 = ~n12202 ;
  assign n12203 = x[32] & n30065 ;
  assign n12204 = n28658 & n12202 ;
  assign n12205 = n12203 | n12204 ;
  assign n12206 = n12198 | n12205 ;
  assign n12207 = n12198 & n12205 ;
  assign n30066 = ~n12207 ;
  assign n12854 = n12206 & n30066 ;
  assign n30067 = ~n12496 ;
  assign n12855 = n30067 & n12854 ;
  assign n30068 = ~n12854 ;
  assign n13064 = n12496 & n30068 ;
  assign n13065 = n12855 | n13064 ;
  assign n4636 = n1720 & n4632 ;
  assign n4553 = x[86] & n4514 ;
  assign n4612 = x[87] & n4572 ;
  assign n13066 = n4553 | n4612 ;
  assign n13067 = x[88] & n4504 ;
  assign n13068 = n13066 | n13067 ;
  assign n13069 = n4636 | n13068 ;
  assign n30069 = ~n13069 ;
  assign n13070 = x[29] & n30069 ;
  assign n13071 = n28483 & n13069 ;
  assign n13072 = n13070 | n13071 ;
  assign n13073 = n13065 | n13072 ;
  assign n13074 = n13065 & n13072 ;
  assign n30070 = ~n13074 ;
  assign n13415 = n13073 & n30070 ;
  assign n30071 = ~n13414 ;
  assign n13416 = n30071 & n13415 ;
  assign n30072 = ~n13415 ;
  assign n13747 = n13414 & n30072 ;
  assign n13748 = n13416 | n13747 ;
  assign n30073 = ~n13746 ;
  assign n14203 = n30073 & n13748 ;
  assign n30074 = ~n13748 ;
  assign n14204 = n13746 & n30074 ;
  assign n14205 = n14203 | n14204 ;
  assign n14206 = n14202 | n14205 ;
  assign n14207 = n14202 & n14205 ;
  assign n30075 = ~n14207 ;
  assign n14644 = n14206 & n30075 ;
  assign n5322 = n2410 & n5302 ;
  assign n5260 = x[92] & n5240 ;
  assign n6239 = x[93] & n6179 ;
  assign n14645 = n5260 | n6239 ;
  assign n14646 = x[94] & n5238 ;
  assign n14647 = n14645 | n14646 ;
  assign n14648 = n5322 | n14647 ;
  assign n30076 = ~n14648 ;
  assign n14649 = x[23] & n30076 ;
  assign n14650 = n28221 & n14648 ;
  assign n14651 = n14649 | n14650 ;
  assign n14652 = n14644 | n14651 ;
  assign n14653 = n14644 & n14651 ;
  assign n30077 = ~n14653 ;
  assign n15542 = n14652 & n30077 ;
  assign n30078 = ~n15144 ;
  assign n15544 = n30078 & n15542 ;
  assign n30079 = ~n15542 ;
  assign n15654 = n15144 & n30079 ;
  assign n15655 = n15544 | n15654 ;
  assign n30080 = ~n15653 ;
  assign n16205 = n30080 & n15655 ;
  assign n30081 = ~n15655 ;
  assign n16511 = n15653 & n30081 ;
  assign n16512 = n16205 | n16511 ;
  assign n16513 = n16510 | n16512 ;
  assign n16514 = n16510 & n16512 ;
  assign n30082 = ~n16514 ;
  assign n16644 = n16513 & n30082 ;
  assign n8760 = n2466 & n8706 ;
  assign n8702 = x[98] & n8645 ;
  assign n9875 = x[99] & n9278 ;
  assign n16645 = n8702 | n9875 ;
  assign n16646 = x[100] & n8643 ;
  assign n16647 = n16645 | n16646 ;
  assign n16648 = n8760 | n16647 ;
  assign n30083 = ~n16648 ;
  assign n16649 = x[17] & n30083 ;
  assign n16650 = n28039 & n16648 ;
  assign n16651 = n16649 | n16650 ;
  assign n16652 = n16644 & n16651 ;
  assign n17169 = n16644 | n16651 ;
  assign n30084 = ~n16652 ;
  assign n17498 = n30084 & n17169 ;
  assign n17499 = n17497 & n17498 ;
  assign n17599 = n17497 | n17498 ;
  assign n30085 = ~n17499 ;
  assign n17600 = n30085 & n17599 ;
  assign n10583 = n2626 & n10542 ;
  assign n10533 = x[101] & n10481 ;
  assign n11881 = x[102] & n11232 ;
  assign n17601 = n10533 | n11881 ;
  assign n17602 = x[103] & n10479 ;
  assign n17603 = n17601 | n17602 ;
  assign n17604 = n10583 | n17603 ;
  assign n30086 = ~n17604 ;
  assign n17605 = x[14] & n30086 ;
  assign n17606 = n27956 & n17604 ;
  assign n17607 = n17605 | n17606 ;
  assign n30087 = ~n17607 ;
  assign n17608 = n17600 & n30087 ;
  assign n30088 = ~n17600 ;
  assign n18690 = n30088 & n17607 ;
  assign n18691 = n17608 | n18690 ;
  assign n17495 = n17450 | n17493 ;
  assign n30089 = ~n17496 ;
  assign n17623 = n17495 & n30089 ;
  assign n18692 = n17620 & n17623 ;
  assign n18761 = n17640 | n18760 ;
  assign n18762 = n18693 & n18761 ;
  assign n18763 = n18692 | n18762 ;
  assign n18764 = n18691 | n18763 ;
  assign n18766 = n18691 & n18763 ;
  assign n30090 = ~n18766 ;
  assign n18833 = n18764 & n30090 ;
  assign n12703 = n3223 & n12695 ;
  assign n12682 = x[104] & n12633 ;
  assign n14371 = x[105] & n13533 ;
  assign n18834 = n12682 | n14371 ;
  assign n18835 = x[106] & n12631 ;
  assign n18836 = n18834 | n18835 ;
  assign n18837 = n12703 | n18836 ;
  assign n30091 = ~n18837 ;
  assign n18838 = x[11] & n30091 ;
  assign n18839 = n27892 & n18837 ;
  assign n18840 = n18838 | n18839 ;
  assign n30092 = ~n18840 ;
  assign n18841 = n18833 & n30092 ;
  assign n30093 = ~n18833 ;
  assign n20041 = n30093 & n18840 ;
  assign n20042 = n18841 | n20041 ;
  assign n30094 = ~n17620 ;
  assign n17624 = n30094 & n17623 ;
  assign n30095 = ~n17623 ;
  assign n17625 = n17620 & n30095 ;
  assign n17626 = n17624 | n17625 ;
  assign n18240 = n17626 | n18239 ;
  assign n18241 = n17626 & n18239 ;
  assign n30096 = ~n18241 ;
  assign n18859 = n18240 & n30096 ;
  assign n20043 = n18856 & n18859 ;
  assign n30097 = ~n18870 ;
  assign n18871 = n18863 & n30097 ;
  assign n30098 = ~n18863 ;
  assign n20046 = n30098 & n18870 ;
  assign n20047 = n18871 | n20046 ;
  assign n20103 = n20047 & n20101 ;
  assign n20104 = n18876 | n20103 ;
  assign n20105 = n20044 & n20104 ;
  assign n20106 = n20043 | n20105 ;
  assign n20107 = n20042 | n20106 ;
  assign n20108 = n20042 & n20106 ;
  assign n30099 = ~n20108 ;
  assign n20147 = n20107 & n30099 ;
  assign n30100 = ~n20146 ;
  assign n20148 = n30100 & n20147 ;
  assign n30101 = ~n20147 ;
  assign n20887 = n20146 & n30101 ;
  assign n20888 = n20148 | n20887 ;
  assign n30102 = ~n20888 ;
  assign n20889 = n20886 & n30102 ;
  assign n21098 = n30020 & n20888 ;
  assign n21099 = n20889 | n21098 ;
  assign n18443 = n4442 & n18392 ;
  assign n18387 = x[110] & n18329 ;
  assign n18565 = x[111] & n18514 ;
  assign n21100 = n18387 | n18565 ;
  assign n21101 = x[112] & n18327 ;
  assign n21102 = n21100 | n21101 ;
  assign n21103 = n18443 | n21102 ;
  assign n30103 = ~n21103 ;
  assign n21104 = x[5] & n30103 ;
  assign n21105 = n27813 & n21103 ;
  assign n21106 = n21104 | n21105 ;
  assign n21107 = n21099 & n21106 ;
  assign n22006 = n21099 | n21106 ;
  assign n30104 = ~n21107 ;
  assign n22294 = n30104 & n22006 ;
  assign n22295 = n22293 & n22294 ;
  assign n22318 = n22293 | n22294 ;
  assign n30105 = ~n22295 ;
  assign n22319 = n30105 & n22318 ;
  assign n30106 = ~n22317 ;
  assign n22320 = n30106 & n22319 ;
  assign n30107 = ~n22319 ;
  assign n23051 = n22317 & n30107 ;
  assign n23052 = n22320 | n23051 ;
  assign n23053 = n23050 | n23052 ;
  assign n23054 = n23050 & n23052 ;
  assign n30108 = ~n23054 ;
  assign n180 = n23053 & n30108 ;
  assign n22321 = n22317 & n22319 ;
  assign n23055 = n22321 | n23054 ;
  assign n22296 = n21107 | n22295 ;
  assign n17609 = n17600 & n17607 ;
  assign n17610 = n17600 | n17607 ;
  assign n30109 = ~n17609 ;
  assign n17611 = n30109 & n17610 ;
  assign n30110 = ~n18763 ;
  assign n18765 = n17611 & n30110 ;
  assign n30111 = ~n17611 ;
  assign n18843 = n30111 & n18763 ;
  assign n18844 = n18765 | n18843 ;
  assign n18846 = n18840 & n18844 ;
  assign n20109 = n18846 | n20108 ;
  assign n18242 = n17622 | n18241 ;
  assign n18243 = n17611 & n18242 ;
  assign n18244 = n17609 | n18243 ;
  assign n8759 = n2977 & n8706 ;
  assign n8704 = x[99] & n8645 ;
  assign n9854 = x[100] & n9278 ;
  assign n16630 = n8704 | n9854 ;
  assign n16631 = x[101] & n8643 ;
  assign n16632 = n16630 | n16631 ;
  assign n16633 = n8759 | n16632 ;
  assign n30112 = ~n16633 ;
  assign n16634 = x[17] & n30112 ;
  assign n16635 = n28039 & n16633 ;
  assign n16636 = n16634 | n16635 ;
  assign n15656 = n15653 & n15655 ;
  assign n16198 = n15688 & n16197 ;
  assign n16199 = n15689 | n16198 ;
  assign n16200 = n15679 & n16199 ;
  assign n16201 = n15677 | n16200 ;
  assign n16203 = n16201 & n16202 ;
  assign n16204 = n15666 | n16203 ;
  assign n16206 = n15653 | n15655 ;
  assign n30113 = ~n15656 ;
  assign n16207 = n30113 & n16206 ;
  assign n16208 = n16204 & n16207 ;
  assign n16209 = n15656 | n16208 ;
  assign n13749 = n13746 & n13748 ;
  assign n14208 = n13749 | n14207 ;
  assign n1842 = n452 & n1841 ;
  assign n350 = x[90] & n330 ;
  assign n432 = x[91] & n390 ;
  assign n13732 = n350 | n432 ;
  assign n13733 = x[92] & n322 ;
  assign n13734 = n13732 | n13733 ;
  assign n13735 = n1842 | n13734 ;
  assign n30114 = ~n13735 ;
  assign n13736 = x[26] & n30114 ;
  assign n13737 = n28342 & n13735 ;
  assign n13738 = n13736 | n13737 ;
  assign n13417 = n13414 & n13415 ;
  assign n13418 = n13074 | n13417 ;
  assign n4648 = n1453 & n4632 ;
  assign n4552 = x[87] & n4514 ;
  assign n4610 = x[88] & n4572 ;
  assign n13055 = n4552 | n4610 ;
  assign n13056 = x[89] & n4504 ;
  assign n13057 = n13055 | n13056 ;
  assign n13058 = n4648 | n13057 ;
  assign n30115 = ~n13058 ;
  assign n13059 = x[29] & n30115 ;
  assign n13060 = n28483 & n13058 ;
  assign n13061 = n13059 | n13060 ;
  assign n3590 = n1270 & n3574 ;
  assign n3503 = x[78] & n3443 ;
  assign n3525 = x[79] & n3508 ;
  assign n10842 = n3503 | n3525 ;
  assign n10843 = x[80] & n3439 ;
  assign n10844 = n10842 | n10843 ;
  assign n10845 = n3590 | n10844 ;
  assign n30116 = ~n10845 ;
  assign n10846 = x[38] & n30116 ;
  assign n10847 = n28996 & n10845 ;
  assign n10848 = n10846 | n10847 ;
  assign n10150 = n10147 & n10149 ;
  assign n10308 = n10150 | n10307 ;
  assign n4796 = n2321 & n4790 ;
  assign n2181 = x[69] & n2179 ;
  assign n2247 = x[70] & n2244 ;
  assign n8980 = n2181 | n2247 ;
  assign n8981 = x[71] & n2175 ;
  assign n8982 = n8980 | n8981 ;
  assign n8983 = n4796 | n8982 ;
  assign n30117 = ~n8983 ;
  assign n8984 = x[47] & n30117 ;
  assign n8985 = n29621 & n8983 ;
  assign n8986 = n8984 | n8985 ;
  assign n8427 = n8418 & n8425 ;
  assign n8428 = n8416 | n8427 ;
  assign n6420 = n2007 & n6408 ;
  assign n1908 = x[66] & n1866 ;
  assign n1951 = x[67] & n1931 ;
  assign n8386 = n1908 | n1951 ;
  assign n8387 = x[68] & n1862 ;
  assign n8388 = n8386 | n8387 ;
  assign n8389 = n6420 | n8388 ;
  assign n8390 = x[50] | n8389 ;
  assign n8391 = x[50] & n8389 ;
  assign n30118 = ~n8391 ;
  assign n8392 = n8390 & n30118 ;
  assign n30119 = ~n7914 ;
  assign n7915 = x[53] & n30119 ;
  assign n27688 = x[52] & x[53] ;
  assign n1545 = x[52] | x[53] ;
  assign n30120 = ~n27688 ;
  assign n1546 = n30120 & n1545 ;
  assign n1690 = n1544 & n1546 ;
  assign n6447 = n1690 & n6437 ;
  assign n30121 = ~n1546 ;
  assign n1547 = n1544 & n30121 ;
  assign n7916 = x[65] & n1547 ;
  assign n27689 = x[51] & x[52] ;
  assign n1548 = x[51] | x[52] ;
  assign n30122 = ~n27689 ;
  assign n1549 = n30122 & n1548 ;
  assign n30123 = ~n1544 ;
  assign n1616 = n30123 & n1549 ;
  assign n7917 = x[64] & n1616 ;
  assign n7918 = n7916 | n7917 ;
  assign n7919 = n6447 | n7918 ;
  assign n30124 = ~n7919 ;
  assign n7920 = x[53] & n30124 ;
  assign n30125 = ~x[53] ;
  assign n7921 = n30125 & n7919 ;
  assign n7922 = n7920 | n7921 ;
  assign n30126 = ~n7922 ;
  assign n7923 = n7915 & n30126 ;
  assign n30127 = ~n7915 ;
  assign n8393 = n30127 & n7922 ;
  assign n8394 = n7923 | n8393 ;
  assign n8395 = n8392 & n8394 ;
  assign n8429 = n8392 | n8394 ;
  assign n30128 = ~n8395 ;
  assign n8430 = n30128 & n8429 ;
  assign n30129 = ~n8428 ;
  assign n8431 = n30129 & n8430 ;
  assign n30130 = ~n8430 ;
  assign n8987 = n8428 & n30130 ;
  assign n8988 = n8431 | n8987 ;
  assign n30131 = ~n8986 ;
  assign n8989 = n30131 & n8988 ;
  assign n30132 = ~n8988 ;
  assign n8991 = n8986 & n30132 ;
  assign n8992 = n8989 | n8991 ;
  assign n9070 = n9004 & n9068 ;
  assign n9071 = n9002 | n9070 ;
  assign n30133 = ~n9071 ;
  assign n9072 = n8992 & n30133 ;
  assign n30134 = ~n8992 ;
  assign n9479 = n30134 & n9071 ;
  assign n9480 = n9072 | n9479 ;
  assign n2727 = n2635 & n2722 ;
  assign n2505 = x[72] & n2492 ;
  assign n2582 = x[73] & n2557 ;
  assign n9481 = n2505 | n2582 ;
  assign n9482 = x[74] & n2488 ;
  assign n9483 = n9481 | n9482 ;
  assign n9484 = n2727 | n9483 ;
  assign n30135 = ~n9484 ;
  assign n9485 = x[44] & n30135 ;
  assign n9486 = n29400 & n9484 ;
  assign n9487 = n9485 | n9486 ;
  assign n9615 = n9480 | n9487 ;
  assign n9488 = n9480 & n9487 ;
  assign n9613 = n9610 & n9611 ;
  assign n9614 = n9499 | n9613 ;
  assign n9617 = n9614 & n9615 ;
  assign n9618 = n9488 | n9617 ;
  assign n30136 = ~n9618 ;
  assign n10127 = n9615 & n30136 ;
  assign n30137 = ~n9488 ;
  assign n9616 = n30137 & n9615 ;
  assign n30138 = ~n9616 ;
  assign n10131 = n9614 & n30138 ;
  assign n10132 = n10127 | n10131 ;
  assign n3168 = n1775 & n3162 ;
  assign n3033 = x[75] & n3031 ;
  assign n3117 = x[76] & n3096 ;
  assign n10133 = n3033 | n3117 ;
  assign n10134 = x[77] & n3027 ;
  assign n10135 = n10133 | n10134 ;
  assign n10136 = n3168 | n10135 ;
  assign n30139 = ~n10136 ;
  assign n10137 = x[41] & n30139 ;
  assign n10138 = n29184 & n10136 ;
  assign n10139 = n10137 | n10138 ;
  assign n10140 = n10132 & n10139 ;
  assign n10309 = n10132 | n10139 ;
  assign n30140 = ~n10140 ;
  assign n10310 = n30140 & n10309 ;
  assign n10311 = n10308 & n10310 ;
  assign n10849 = n10308 | n10310 ;
  assign n30141 = ~n10311 ;
  assign n10850 = n30141 & n10849 ;
  assign n30142 = ~n10848 ;
  assign n10851 = n30142 & n10850 ;
  assign n30143 = ~n10850 ;
  assign n10853 = n10848 & n30143 ;
  assign n10854 = n10851 | n10853 ;
  assign n11073 = n10866 | n11072 ;
  assign n11074 = n10854 | n11073 ;
  assign n11075 = n10854 & n11073 ;
  assign n30144 = ~n11075 ;
  assign n11412 = n11074 & n30144 ;
  assign n4082 = n1057 & n4041 ;
  assign n3921 = x[81] & n3910 ;
  assign n4013 = x[82] & n3975 ;
  assign n11413 = n3921 | n4013 ;
  assign n11414 = x[83] & n3906 ;
  assign n11415 = n11413 | n11414 ;
  assign n11416 = n4082 | n11415 ;
  assign n30145 = ~n11416 ;
  assign n11417 = x[35] & n30145 ;
  assign n11418 = n28822 & n11416 ;
  assign n11419 = n11417 | n11418 ;
  assign n11680 = n11412 | n11419 ;
  assign n11420 = n11412 & n11419 ;
  assign n12180 = n11676 & n12178 ;
  assign n12181 = n11430 | n12180 ;
  assign n12182 = n11680 & n12181 ;
  assign n12183 = n11420 | n12182 ;
  assign n30146 = ~n12183 ;
  assign n12184 = n11680 & n30146 ;
  assign n11653 = n11649 & n11652 ;
  assign n11654 = n11511 | n11653 ;
  assign n11656 = n11498 | n11500 ;
  assign n30147 = ~n11501 ;
  assign n11657 = n30147 & n11656 ;
  assign n11658 = n11654 & n11657 ;
  assign n11659 = n11501 | n11658 ;
  assign n11660 = n11490 & n11659 ;
  assign n11661 = n11491 | n11660 ;
  assign n11663 = n11471 | n11473 ;
  assign n30148 = ~n11474 ;
  assign n11664 = n30148 & n11663 ;
  assign n11665 = n11661 & n11664 ;
  assign n11666 = n11474 | n11665 ;
  assign n11667 = n11463 & n11666 ;
  assign n11668 = n11464 | n11667 ;
  assign n11669 = n11452 & n11668 ;
  assign n11670 = n11449 | n11669 ;
  assign n11674 = n11670 & n11673 ;
  assign n11675 = n11439 | n11674 ;
  assign n11678 = n11675 & n11677 ;
  assign n11679 = n11430 | n11678 ;
  assign n30149 = ~n11420 ;
  assign n12141 = n30149 & n11680 ;
  assign n30150 = ~n12141 ;
  assign n12185 = n11679 & n30150 ;
  assign n12186 = n12184 | n12185 ;
  assign n1214 = n779 & n1213 ;
  assign n707 = x[84] & n663 ;
  assign n756 = x[85] & n720 ;
  assign n12187 = n707 | n756 ;
  assign n12188 = x[86] & n652 ;
  assign n12189 = n12187 | n12188 ;
  assign n12190 = n1214 | n12189 ;
  assign n30151 = ~n12190 ;
  assign n12191 = x[32] & n30151 ;
  assign n12192 = n28658 & n12190 ;
  assign n12193 = n12191 | n12192 ;
  assign n12194 = n12186 | n12193 ;
  assign n12195 = n12186 & n12193 ;
  assign n30152 = ~n12195 ;
  assign n12196 = n12194 & n30152 ;
  assign n12899 = n12221 | n12898 ;
  assign n12900 = n12854 & n12899 ;
  assign n12901 = n12207 | n12900 ;
  assign n12903 = n12196 | n12901 ;
  assign n12904 = n12196 & n12901 ;
  assign n30153 = ~n12904 ;
  assign n13419 = n12903 & n30153 ;
  assign n30154 = ~n13061 ;
  assign n13420 = n30154 & n13419 ;
  assign n30155 = ~n13419 ;
  assign n13421 = n13061 & n30155 ;
  assign n13422 = n13420 | n13421 ;
  assign n30156 = ~n13422 ;
  assign n13658 = n13418 & n30156 ;
  assign n30157 = ~n13418 ;
  assign n14209 = n30157 & n13422 ;
  assign n14210 = n13658 | n14209 ;
  assign n14211 = n13738 | n14210 ;
  assign n14212 = n13738 & n14210 ;
  assign n30158 = ~n14212 ;
  assign n14213 = n14211 & n30158 ;
  assign n14214 = n14208 & n14213 ;
  assign n14631 = n14208 | n14213 ;
  assign n30159 = ~n14214 ;
  assign n14632 = n30159 & n14631 ;
  assign n5324 = n2152 & n5302 ;
  assign n5243 = x[93] & n5240 ;
  assign n6243 = x[94] & n6179 ;
  assign n14633 = n5243 | n6243 ;
  assign n14634 = x[95] & n5238 ;
  assign n14635 = n14633 | n14634 ;
  assign n14636 = n5324 | n14635 ;
  assign n30160 = ~n14636 ;
  assign n14637 = x[23] & n30160 ;
  assign n14638 = n28221 & n14636 ;
  assign n14639 = n14637 | n14638 ;
  assign n14641 = n14632 & n14639 ;
  assign n14642 = n14632 | n14639 ;
  assign n30161 = ~n14641 ;
  assign n14643 = n30161 & n14642 ;
  assign n15136 = n14670 & n15134 ;
  assign n15536 = n14670 | n15134 ;
  assign n30162 = ~n15136 ;
  assign n15537 = n30162 & n15536 ;
  assign n15538 = n15534 & n15537 ;
  assign n15539 = n14673 | n15538 ;
  assign n15540 = n15141 & n15539 ;
  assign n15541 = n14663 | n15540 ;
  assign n15543 = n15541 & n15542 ;
  assign n15545 = n14653 | n15543 ;
  assign n30163 = ~n15545 ;
  assign n15546 = n14643 & n30163 ;
  assign n30164 = ~n14643 ;
  assign n15632 = n30164 & n15545 ;
  assign n15633 = n15546 | n15632 ;
  assign n7205 = n2841 & n7162 ;
  assign n7119 = x[96] & n7100 ;
  assign n7705 = x[97] & n7647 ;
  assign n15634 = n7119 | n7705 ;
  assign n15635 = x[98] & n7098 ;
  assign n15636 = n15634 | n15635 ;
  assign n15637 = n7205 | n15636 ;
  assign n30165 = ~n15637 ;
  assign n15638 = x[20] & n30165 ;
  assign n15639 = n28114 & n15637 ;
  assign n15640 = n15638 | n15639 ;
  assign n15641 = n15633 | n15640 ;
  assign n15642 = n15633 & n15640 ;
  assign n30166 = ~n15642 ;
  assign n16398 = n15641 & n30166 ;
  assign n30167 = ~n16209 ;
  assign n16399 = n30167 & n16398 ;
  assign n30168 = ~n16398 ;
  assign n16639 = n16209 & n30168 ;
  assign n16640 = n16399 | n16639 ;
  assign n16641 = n16636 | n16640 ;
  assign n16642 = n16636 & n16640 ;
  assign n30169 = ~n16642 ;
  assign n16643 = n16641 & n30169 ;
  assign n17500 = n16652 | n17499 ;
  assign n30170 = ~n17500 ;
  assign n17501 = n16643 & n30170 ;
  assign n30171 = ~n16643 ;
  assign n17584 = n30171 & n17500 ;
  assign n17585 = n17501 | n17584 ;
  assign n10577 = n3001 & n10542 ;
  assign n10540 = x[102] & n10481 ;
  assign n11883 = x[103] & n11232 ;
  assign n17586 = n10540 | n11883 ;
  assign n17587 = x[104] & n10479 ;
  assign n17588 = n17586 | n17587 ;
  assign n17589 = n10577 | n17588 ;
  assign n30172 = ~n17589 ;
  assign n17590 = x[14] & n30172 ;
  assign n17591 = n27956 & n17589 ;
  assign n17592 = n17590 | n17591 ;
  assign n17593 = n17585 | n17592 ;
  assign n17594 = n17585 & n17592 ;
  assign n30173 = ~n17594 ;
  assign n18688 = n17593 & n30173 ;
  assign n30174 = ~n18244 ;
  assign n18689 = n30174 & n18688 ;
  assign n30175 = ~n18688 ;
  assign n18823 = n18244 & n30175 ;
  assign n18824 = n18689 | n18823 ;
  assign n12753 = n3199 & n12695 ;
  assign n12686 = x[105] & n12633 ;
  assign n14391 = x[106] & n13533 ;
  assign n18825 = n12686 | n14391 ;
  assign n18826 = x[107] & n12631 ;
  assign n18827 = n18825 | n18826 ;
  assign n18828 = n12753 | n18827 ;
  assign n30176 = ~n18828 ;
  assign n18829 = x[11] & n30176 ;
  assign n18830 = n27892 & n18828 ;
  assign n18831 = n18829 | n18830 ;
  assign n19542 = n18824 | n18831 ;
  assign n30177 = ~n14639 ;
  assign n14640 = n14632 & n30177 ;
  assign n30178 = ~n14632 ;
  assign n15518 = n30178 & n14639 ;
  assign n15519 = n14640 | n15518 ;
  assign n15547 = n15519 | n15545 ;
  assign n15548 = n15519 & n15545 ;
  assign n30179 = ~n15548 ;
  assign n15643 = n15547 & n30179 ;
  assign n30180 = ~n15640 ;
  assign n15644 = n30180 & n15643 ;
  assign n30181 = ~n15643 ;
  assign n15645 = n15640 & n30181 ;
  assign n15646 = n15644 | n15645 ;
  assign n16210 = n15646 | n16209 ;
  assign n16211 = n15646 & n16209 ;
  assign n30182 = ~n16211 ;
  assign n16629 = n16210 & n30182 ;
  assign n30183 = ~n16636 ;
  assign n16637 = n16629 & n30183 ;
  assign n30184 = ~n16629 ;
  assign n17447 = n30184 & n16636 ;
  assign n17448 = n16637 | n17447 ;
  assign n17502 = n17448 | n17500 ;
  assign n17503 = n17448 & n17500 ;
  assign n30185 = ~n17503 ;
  assign n17595 = n17502 & n30185 ;
  assign n30186 = ~n17592 ;
  assign n17596 = n30186 & n17595 ;
  assign n30187 = ~n17595 ;
  assign n17597 = n17592 & n30187 ;
  assign n17598 = n17596 | n17597 ;
  assign n18245 = n17598 | n18244 ;
  assign n18246 = n17598 & n18244 ;
  assign n30188 = ~n18246 ;
  assign n20039 = n18245 & n30188 ;
  assign n20040 = n18831 & n20039 ;
  assign n30189 = ~n20040 ;
  assign n20125 = n19542 & n30189 ;
  assign n30190 = ~n20125 ;
  assign n20126 = n20109 & n30190 ;
  assign n18832 = n18824 & n18831 ;
  assign n18842 = n18833 & n18840 ;
  assign n18845 = n18840 | n18844 ;
  assign n30191 = ~n18846 ;
  assign n18847 = n18845 & n30191 ;
  assign n30192 = ~n18856 ;
  assign n18860 = n30192 & n18859 ;
  assign n30193 = ~n18859 ;
  assign n18861 = n18856 & n30193 ;
  assign n18862 = n18860 | n18861 ;
  assign n19538 = n18862 & n19537 ;
  assign n19539 = n18858 | n19538 ;
  assign n19540 = n18847 & n19539 ;
  assign n19541 = n18842 | n19540 ;
  assign n19543 = n19541 & n19542 ;
  assign n19544 = n18832 | n19543 ;
  assign n30194 = ~n19544 ;
  assign n20127 = n19542 & n30194 ;
  assign n20128 = n20126 | n20127 ;
  assign n15322 = n3615 & n15308 ;
  assign n15258 = x[108] & n15246 ;
  assign n17325 = x[109] & n16288 ;
  assign n20129 = n15258 | n17325 ;
  assign n20130 = x[110] & n15244 ;
  assign n20131 = n20129 | n20130 ;
  assign n20132 = n15322 | n20131 ;
  assign n30195 = ~n20132 ;
  assign n20133 = x[8] & n30195 ;
  assign n20134 = n27845 & n20132 ;
  assign n20135 = n20133 | n20134 ;
  assign n30196 = ~n20135 ;
  assign n20136 = n20128 & n30196 ;
  assign n30197 = ~n20128 ;
  assign n20138 = n30197 & n20135 ;
  assign n20139 = n20136 | n20138 ;
  assign n20149 = n20146 & n20147 ;
  assign n20890 = n20886 & n20888 ;
  assign n20891 = n20149 | n20890 ;
  assign n20892 = n20139 | n20891 ;
  assign n20893 = n20139 & n20891 ;
  assign n30198 = ~n20893 ;
  assign n21088 = n20892 & n30198 ;
  assign n18441 = n4087 & n18392 ;
  assign n18375 = x[111] & n18329 ;
  assign n18562 = x[112] & n18514 ;
  assign n21089 = n18375 | n18562 ;
  assign n21090 = x[113] & n18327 ;
  assign n21091 = n21089 | n21090 ;
  assign n21092 = n18441 | n21091 ;
  assign n30199 = ~n21092 ;
  assign n21093 = x[5] & n30199 ;
  assign n21094 = n27813 & n21092 ;
  assign n21095 = n21093 | n21094 ;
  assign n30200 = ~n21095 ;
  assign n21096 = n21088 & n30200 ;
  assign n30201 = ~n21088 ;
  assign n22297 = n30201 & n21095 ;
  assign n22298 = n21096 | n22297 ;
  assign n22299 = n22296 | n22298 ;
  assign n22300 = n22296 & n22298 ;
  assign n30202 = ~n22300 ;
  assign n22301 = n22299 & n30202 ;
  assign n609 = n607 & n608 ;
  assign n610 = n27592 | n609 ;
  assign n24199 = x[115] & x[116] ;
  assign n611 = x[115] | x[116] ;
  assign n30203 = ~n24199 ;
  assign n4699 = n30203 & n611 ;
  assign n4700 = n610 & n4699 ;
  assign n4701 = n610 | n4699 ;
  assign n30204 = ~n4700 ;
  assign n4702 = n30204 & n4701 ;
  assign n19694 = n4702 & n19656 ;
  assign n19752 = x[114] & n19723 ;
  assign n19866 = x[115] & n19829 ;
  assign n22302 = n19752 | n19866 ;
  assign n22303 = x[116] & n19655 ;
  assign n22304 = n22302 | n22303 ;
  assign n22305 = n19694 | n22304 ;
  assign n30205 = ~n22305 ;
  assign n22306 = x[2] & n30205 ;
  assign n22307 = n27790 & n22305 ;
  assign n22308 = n22306 | n22307 ;
  assign n22309 = n22301 | n22308 ;
  assign n22310 = n22301 & n22308 ;
  assign n30206 = ~n22310 ;
  assign n23056 = n22309 & n30206 ;
  assign n23057 = n23055 & n23056 ;
  assign n27699 = n23055 | n23056 ;
  assign n30207 = ~n23057 ;
  assign n181 = n30207 & n27699 ;
  assign n23058 = n22310 | n23057 ;
  assign n21097 = n21088 & n21095 ;
  assign n23059 = n21097 | n22300 ;
  assign n8750 = n2867 & n8706 ;
  assign n8698 = x[100] & n8645 ;
  assign n9876 = x[101] & n9278 ;
  assign n16616 = n8698 | n9876 ;
  assign n16617 = x[102] & n8643 ;
  assign n16618 = n16616 | n16617 ;
  assign n16619 = n8750 | n16618 ;
  assign n30208 = ~n16619 ;
  assign n16620 = x[17] & n30208 ;
  assign n16621 = n28039 & n16619 ;
  assign n16622 = n16620 | n16621 ;
  assign n7183 = n2313 & n7162 ;
  assign n7123 = x[97] & n7100 ;
  assign n7703 = x[98] & n7647 ;
  assign n15619 = n7123 | n7703 ;
  assign n15620 = x[99] & n7098 ;
  assign n15621 = n15619 | n15620 ;
  assign n15622 = n7183 | n15621 ;
  assign n30209 = ~n15622 ;
  assign n15623 = x[20] & n30209 ;
  assign n15624 = n28114 & n15622 ;
  assign n15625 = n15623 | n15624 ;
  assign n15549 = n14641 | n15548 ;
  assign n5326 = n2000 & n5302 ;
  assign n5261 = x[94] & n5240 ;
  assign n6254 = x[95] & n6179 ;
  assign n14621 = n5261 | n6254 ;
  assign n14622 = x[96] & n5238 ;
  assign n14623 = n14621 | n14622 ;
  assign n14624 = n5326 | n14623 ;
  assign n30210 = ~n14624 ;
  assign n14625 = x[23] & n30210 ;
  assign n14626 = n28221 & n14624 ;
  assign n14627 = n14625 | n14626 ;
  assign n13423 = n13418 | n13422 ;
  assign n13424 = n13418 & n13422 ;
  assign n30211 = ~n13424 ;
  assign n13731 = n13423 & n30211 ;
  assign n13739 = n13731 & n13738 ;
  assign n14215 = n13739 | n14214 ;
  assign n1686 = n452 & n1685 ;
  assign n353 = x[91] & n330 ;
  assign n430 = x[92] & n390 ;
  assign n13721 = n353 | n430 ;
  assign n13722 = x[93] & n322 ;
  assign n13723 = n13721 | n13722 ;
  assign n13724 = n1686 | n13723 ;
  assign n30212 = ~n13724 ;
  assign n13725 = x[26] & n30212 ;
  assign n13726 = n28342 & n13724 ;
  assign n13727 = n13725 | n13726 ;
  assign n30213 = ~n12901 ;
  assign n12902 = n12196 & n30213 ;
  assign n30214 = ~n12196 ;
  assign n13053 = n30214 & n12901 ;
  assign n13054 = n12902 | n13053 ;
  assign n13063 = n13054 & n13061 ;
  assign n13425 = n13063 | n13424 ;
  assign n1524 = n779 & n1522 ;
  assign n705 = x[85] & n663 ;
  assign n729 = x[86] & n720 ;
  assign n12131 = n705 | n729 ;
  assign n12132 = x[87] & n652 ;
  assign n12133 = n12131 | n12132 ;
  assign n12134 = n1524 | n12133 ;
  assign n30215 = ~n12134 ;
  assign n12135 = x[32] & n30215 ;
  assign n12136 = n28658 & n12134 ;
  assign n12137 = n12135 | n12136 ;
  assign n11681 = n11679 & n11680 ;
  assign n11682 = n11420 | n11681 ;
  assign n10852 = n10848 & n10850 ;
  assign n11076 = n10852 | n11075 ;
  assign n3581 = n1029 & n3574 ;
  assign n3465 = x[79] & n3443 ;
  assign n3542 = x[80] & n3508 ;
  assign n10832 = n3465 | n3542 ;
  assign n10833 = x[81] & n3439 ;
  assign n10834 = n10832 | n10833 ;
  assign n10835 = n3581 | n10834 ;
  assign n30216 = ~n10835 ;
  assign n10836 = x[38] & n30216 ;
  assign n10837 = n28996 & n10835 ;
  assign n10838 = n10836 | n10837 ;
  assign n10312 = n10140 | n10311 ;
  assign n3163 = n2084 & n3162 ;
  assign n3064 = x[76] & n3031 ;
  assign n3119 = x[77] & n3096 ;
  assign n10119 = n3064 | n3119 ;
  assign n10120 = x[78] & n3027 ;
  assign n10121 = n10119 | n10120 ;
  assign n10122 = n3163 | n10121 ;
  assign n30217 = ~n10122 ;
  assign n10123 = x[41] & n30217 ;
  assign n10124 = n29184 & n10122 ;
  assign n10125 = n10123 | n10124 ;
  assign n3294 = n2635 & n3289 ;
  assign n2521 = x[73] & n2492 ;
  assign n2583 = x[74] & n2557 ;
  assign n9468 = n2521 | n2583 ;
  assign n9469 = x[75] & n2488 ;
  assign n9470 = n9468 | n9469 ;
  assign n9471 = n3294 | n9470 ;
  assign n30218 = ~n9471 ;
  assign n9472 = x[44] & n30218 ;
  assign n9473 = n29400 & n9471 ;
  assign n9474 = n9472 | n9473 ;
  assign n8990 = n8986 & n8988 ;
  assign n9073 = n8992 & n9071 ;
  assign n9074 = n8990 | n9073 ;
  assign n8432 = n8428 & n8430 ;
  assign n8433 = n8395 | n8432 ;
  assign n7924 = n7915 & n7922 ;
  assign n6475 = n1690 & n6466 ;
  assign n1550 = n30123 & n1546 ;
  assign n30219 = ~n1549 ;
  assign n1551 = n30219 & n1550 ;
  assign n1575 = x[64] & n1551 ;
  assign n1623 = x[65] & n1616 ;
  assign n7925 = n1575 | n1623 ;
  assign n7926 = x[66] & n1547 ;
  assign n7927 = n7925 | n7926 ;
  assign n7928 = n6475 | n7927 ;
  assign n30220 = ~n7928 ;
  assign n7929 = x[53] & n30220 ;
  assign n7930 = n30125 & n7928 ;
  assign n7931 = n7929 | n7930 ;
  assign n30221 = ~n7931 ;
  assign n7932 = n7924 & n30221 ;
  assign n30222 = ~n7924 ;
  assign n8376 = n30222 & n7931 ;
  assign n8377 = n7932 | n8376 ;
  assign n6385 = n2007 & n6379 ;
  assign n1876 = x[67] & n1866 ;
  assign n1953 = x[68] & n1931 ;
  assign n8378 = n1876 | n1953 ;
  assign n8379 = x[69] & n1862 ;
  assign n8380 = n8378 | n8379 ;
  assign n8381 = n6385 | n8380 ;
  assign n30223 = ~n8381 ;
  assign n8382 = x[50] & n30223 ;
  assign n8383 = n29865 & n8381 ;
  assign n8384 = n8382 | n8383 ;
  assign n8385 = n8377 & n8384 ;
  assign n8434 = n8377 | n8384 ;
  assign n30224 = ~n8385 ;
  assign n8435 = n30224 & n8434 ;
  assign n30225 = ~n8435 ;
  assign n8969 = n8433 & n30225 ;
  assign n8436 = n8433 & n8434 ;
  assign n8437 = n8385 | n8436 ;
  assign n30226 = ~n8437 ;
  assign n8970 = n8434 & n30226 ;
  assign n8971 = n8969 | n8970 ;
  assign n3709 = n2321 & n3701 ;
  assign n2193 = x[70] & n2179 ;
  assign n2265 = x[71] & n2244 ;
  assign n8972 = n2193 | n2265 ;
  assign n8973 = x[72] & n2175 ;
  assign n8974 = n8972 | n8973 ;
  assign n8975 = n3709 | n8974 ;
  assign n30227 = ~n8975 ;
  assign n8976 = x[47] & n30227 ;
  assign n8977 = n29621 & n8975 ;
  assign n8978 = n8976 | n8977 ;
  assign n8979 = n8971 | n8978 ;
  assign n9075 = n8971 & n8978 ;
  assign n30228 = ~n9075 ;
  assign n9076 = n8979 & n30228 ;
  assign n9077 = n9074 & n9076 ;
  assign n9475 = n9074 | n9076 ;
  assign n30229 = ~n9077 ;
  assign n9476 = n30229 & n9475 ;
  assign n30230 = ~n9474 ;
  assign n9477 = n30230 & n9476 ;
  assign n30231 = ~n9476 ;
  assign n9619 = n9474 & n30231 ;
  assign n9620 = n9477 | n9619 ;
  assign n9621 = n9618 & n9620 ;
  assign n10313 = n9618 | n9620 ;
  assign n30232 = ~n9621 ;
  assign n10314 = n30232 & n10313 ;
  assign n30233 = ~n10125 ;
  assign n10315 = n30233 & n10314 ;
  assign n30234 = ~n10314 ;
  assign n10317 = n10125 & n30234 ;
  assign n10318 = n10315 | n10317 ;
  assign n10319 = n10312 | n10318 ;
  assign n10320 = n10312 & n10318 ;
  assign n30235 = ~n10320 ;
  assign n10839 = n10319 & n30235 ;
  assign n30236 = ~n10838 ;
  assign n10840 = n30236 & n10839 ;
  assign n30237 = ~n10839 ;
  assign n11077 = n10838 & n30237 ;
  assign n11078 = n10840 | n11077 ;
  assign n11079 = n11076 & n11078 ;
  assign n11401 = n11076 | n11078 ;
  assign n30238 = ~n11079 ;
  assign n11402 = n30238 & n11401 ;
  assign n4071 = n1293 & n4041 ;
  assign n3932 = x[82] & n3910 ;
  assign n3997 = x[83] & n3975 ;
  assign n11403 = n3932 | n3997 ;
  assign n11404 = x[84] & n3906 ;
  assign n11405 = n11403 | n11404 ;
  assign n11406 = n4071 | n11405 ;
  assign n30239 = ~n11406 ;
  assign n11407 = x[35] & n30239 ;
  assign n11408 = n28822 & n11406 ;
  assign n11409 = n11407 | n11408 ;
  assign n30240 = ~n11409 ;
  assign n11410 = n11402 & n30240 ;
  assign n30241 = ~n11402 ;
  assign n11683 = n30241 & n11409 ;
  assign n11684 = n11410 | n11683 ;
  assign n30242 = ~n11684 ;
  assign n11685 = n11682 & n30242 ;
  assign n30243 = ~n11682 ;
  assign n12138 = n30243 & n11684 ;
  assign n12139 = n11685 | n12138 ;
  assign n30244 = ~n12137 ;
  assign n12501 = n30244 & n12139 ;
  assign n30245 = ~n12139 ;
  assign n12502 = n12137 & n30245 ;
  assign n12503 = n12501 | n12502 ;
  assign n12905 = n12195 | n12904 ;
  assign n30246 = ~n12503 ;
  assign n12906 = n30246 & n12905 ;
  assign n30247 = ~n12905 ;
  assign n13043 = n12503 & n30247 ;
  assign n13044 = n12906 | n13043 ;
  assign n4649 = n1482 & n4632 ;
  assign n4536 = x[88] & n4514 ;
  assign n4573 = x[89] & n4572 ;
  assign n13045 = n4536 | n4573 ;
  assign n13046 = x[90] & n4504 ;
  assign n13047 = n13045 | n13046 ;
  assign n13048 = n4649 | n13047 ;
  assign n30248 = ~n13048 ;
  assign n13049 = x[29] & n30248 ;
  assign n13050 = n28483 & n13048 ;
  assign n13051 = n13049 | n13050 ;
  assign n13052 = n13044 & n13051 ;
  assign n13426 = n13044 | n13051 ;
  assign n30249 = ~n13052 ;
  assign n13427 = n30249 & n13426 ;
  assign n13428 = n13425 & n13427 ;
  assign n13728 = n13425 | n13427 ;
  assign n30250 = ~n13428 ;
  assign n13729 = n30250 & n13728 ;
  assign n13730 = n13727 & n13729 ;
  assign n14216 = n13727 | n13729 ;
  assign n30251 = ~n13730 ;
  assign n14605 = n30251 & n14216 ;
  assign n30252 = ~n14215 ;
  assign n14607 = n30252 & n14605 ;
  assign n30253 = ~n14605 ;
  assign n14628 = n14215 & n30253 ;
  assign n14629 = n14607 | n14628 ;
  assign n14630 = n14627 & n14629 ;
  assign n15149 = n14627 | n14629 ;
  assign n30254 = ~n14630 ;
  assign n15550 = n30254 & n15149 ;
  assign n15551 = n15549 & n15550 ;
  assign n15626 = n15549 | n15550 ;
  assign n30255 = ~n15551 ;
  assign n15627 = n30255 & n15626 ;
  assign n30256 = ~n15625 ;
  assign n15629 = n30256 & n15627 ;
  assign n30257 = ~n15627 ;
  assign n16395 = n15625 & n30257 ;
  assign n16396 = n15629 | n16395 ;
  assign n16397 = n15640 & n15643 ;
  assign n16515 = n15656 | n16514 ;
  assign n16516 = n16398 & n16515 ;
  assign n16517 = n16397 | n16516 ;
  assign n16519 = n16396 | n16517 ;
  assign n16520 = n16396 & n16517 ;
  assign n30258 = ~n16520 ;
  assign n16625 = n16519 & n30258 ;
  assign n30259 = ~n16622 ;
  assign n16626 = n30259 & n16625 ;
  assign n30260 = ~n16625 ;
  assign n16627 = n16622 & n30260 ;
  assign n16628 = n16626 | n16627 ;
  assign n16638 = n16629 & n16636 ;
  assign n17166 = n16676 | n17165 ;
  assign n17167 = n16665 & n17166 ;
  assign n17168 = n16662 | n17167 ;
  assign n17170 = n17168 & n17169 ;
  assign n17171 = n16652 | n17170 ;
  assign n17172 = n16643 & n17171 ;
  assign n17173 = n16638 | n17172 ;
  assign n17174 = n16628 | n17173 ;
  assign n17175 = n16628 & n17173 ;
  assign n30261 = ~n17175 ;
  assign n17569 = n17174 & n30261 ;
  assign n10601 = n3409 & n10542 ;
  assign n10516 = x[103] & n10481 ;
  assign n11887 = x[104] & n11232 ;
  assign n17570 = n10516 | n11887 ;
  assign n17571 = x[105] & n10479 ;
  assign n17572 = n17570 | n17571 ;
  assign n17573 = n10601 | n17572 ;
  assign n30262 = ~n17573 ;
  assign n17574 = x[14] & n30262 ;
  assign n17575 = n27956 & n17573 ;
  assign n17576 = n17574 | n17575 ;
  assign n30263 = ~n17576 ;
  assign n17577 = n17569 & n30263 ;
  assign n30264 = ~n17569 ;
  assign n18685 = n30264 & n17576 ;
  assign n18686 = n17577 | n18685 ;
  assign n18687 = n17592 & n17595 ;
  assign n18767 = n17609 | n18766 ;
  assign n18768 = n18688 & n18767 ;
  assign n18769 = n18687 | n18768 ;
  assign n18770 = n18686 | n18769 ;
  assign n18771 = n18686 & n18769 ;
  assign n30265 = ~n18771 ;
  assign n18814 = n18770 & n30265 ;
  assign n12739 = n3876 & n12695 ;
  assign n12674 = x[106] & n12633 ;
  assign n14396 = x[107] & n13533 ;
  assign n18815 = n12674 | n14396 ;
  assign n18816 = x[108] & n12631 ;
  assign n18817 = n18815 | n18816 ;
  assign n18818 = n12739 | n18817 ;
  assign n30266 = ~n18818 ;
  assign n18819 = x[11] & n30266 ;
  assign n18820 = n27892 & n18818 ;
  assign n18821 = n18819 | n18820 ;
  assign n19545 = n18814 | n18821 ;
  assign n18822 = n18814 & n18821 ;
  assign n19546 = n19544 & n19545 ;
  assign n19547 = n18822 | n19546 ;
  assign n30267 = ~n19547 ;
  assign n19548 = n19545 & n30267 ;
  assign n30268 = ~n18822 ;
  assign n20038 = n30268 & n19545 ;
  assign n20110 = n18831 | n20039 ;
  assign n20111 = n20109 & n20110 ;
  assign n20112 = n20040 | n20111 ;
  assign n30269 = ~n20038 ;
  assign n20113 = n30269 & n20112 ;
  assign n20114 = n19548 | n20113 ;
  assign n15345 = n4246 & n15308 ;
  assign n15296 = x[109] & n15246 ;
  assign n17320 = x[110] & n16288 ;
  assign n20115 = n15296 | n17320 ;
  assign n20116 = x[111] & n15244 ;
  assign n20117 = n20115 | n20116 ;
  assign n20118 = n15345 | n20117 ;
  assign n30270 = ~n20118 ;
  assign n20119 = x[8] & n30270 ;
  assign n20120 = n27845 & n20118 ;
  assign n20121 = n20119 | n20120 ;
  assign n20122 = n20114 | n20121 ;
  assign n20123 = n20114 & n20121 ;
  assign n30271 = ~n20123 ;
  assign n20124 = n20122 & n30271 ;
  assign n20137 = n20128 & n20135 ;
  assign n20894 = n20137 | n20893 ;
  assign n20895 = n20124 & n20894 ;
  assign n21078 = n20124 | n20894 ;
  assign n30272 = ~n20895 ;
  assign n21079 = n30272 & n21078 ;
  assign n18428 = n4276 & n18392 ;
  assign n18389 = x[112] & n18329 ;
  assign n18539 = x[113] & n18514 ;
  assign n21080 = n18389 | n18539 ;
  assign n21081 = x[114] & n18327 ;
  assign n21082 = n21080 | n21081 ;
  assign n21083 = n18428 | n21082 ;
  assign n30273 = ~n21083 ;
  assign n21084 = x[5] & n30273 ;
  assign n21085 = n27813 & n21083 ;
  assign n21086 = n21084 | n21085 ;
  assign n21087 = n21079 & n21086 ;
  assign n22013 = n21079 | n21086 ;
  assign n30274 = ~n21087 ;
  assign n23060 = n30274 & n22013 ;
  assign n30275 = ~n23060 ;
  assign n23061 = n23059 & n30275 ;
  assign n30276 = ~n21317 ;
  assign n21322 = n30276 & n21321 ;
  assign n30277 = ~n21321 ;
  assign n21323 = n21317 & n30277 ;
  assign n21324 = n21322 | n21323 ;
  assign n22002 = n21324 & n22001 ;
  assign n22003 = n21319 | n22002 ;
  assign n22004 = n21308 & n22003 ;
  assign n22005 = n21306 | n22004 ;
  assign n22007 = n22005 & n22006 ;
  assign n22008 = n21107 | n22007 ;
  assign n22009 = n21088 | n21095 ;
  assign n30278 = ~n21097 ;
  assign n22010 = n30278 & n22009 ;
  assign n22011 = n22008 & n22010 ;
  assign n22012 = n21097 | n22011 ;
  assign n22014 = n22012 & n22013 ;
  assign n22015 = n21087 | n22014 ;
  assign n30279 = ~n22015 ;
  assign n23062 = n22013 & n30279 ;
  assign n23063 = n23061 | n23062 ;
  assign n612 = n610 & n611 ;
  assign n613 = n24199 | n612 ;
  assign n27570 = x[116] & x[117] ;
  assign n614 = x[116] | x[117] ;
  assign n30280 = ~n27570 ;
  assign n794 = n30280 & n614 ;
  assign n30281 = ~n613 ;
  assign n795 = n30281 & n794 ;
  assign n30282 = ~n794 ;
  assign n796 = n613 & n30282 ;
  assign n797 = n795 | n796 ;
  assign n19721 = n797 & n19656 ;
  assign n19787 = x[115] & n19723 ;
  assign n19863 = x[116] & n19829 ;
  assign n23064 = n19787 | n19863 ;
  assign n23065 = x[117] & n19655 ;
  assign n23066 = n23064 | n23065 ;
  assign n23067 = n19721 | n23066 ;
  assign n30283 = ~n23067 ;
  assign n23068 = x[2] & n30283 ;
  assign n23069 = n27790 & n23067 ;
  assign n23070 = n23068 | n23069 ;
  assign n30284 = ~n23070 ;
  assign n23071 = n23063 & n30284 ;
  assign n30285 = ~n23063 ;
  assign n23072 = n30285 & n23070 ;
  assign n23073 = n23071 | n23072 ;
  assign n23074 = n23058 | n23073 ;
  assign n23076 = n23058 & n23073 ;
  assign n30286 = ~n23076 ;
  assign n182 = n23074 & n30286 ;
  assign n23075 = n23063 & n23070 ;
  assign n23077 = n23075 | n23076 ;
  assign n615 = n613 & n614 ;
  assign n616 = n27570 | n615 ;
  assign n24007 = x[117] & x[118] ;
  assign n617 = x[117] | x[118] ;
  assign n30287 = ~n24007 ;
  assign n781 = n30287 & n617 ;
  assign n782 = n616 & n781 ;
  assign n783 = n616 | n781 ;
  assign n30288 = ~n782 ;
  assign n784 = n30288 & n783 ;
  assign n19678 = n784 & n19656 ;
  assign n19780 = x[116] & n19723 ;
  assign n19870 = x[117] & n19829 ;
  assign n22086 = n19780 | n19870 ;
  assign n22087 = x[118] & n19655 ;
  assign n22088 = n22086 | n22087 ;
  assign n22089 = n19678 | n22088 ;
  assign n22090 = x[2] | n22089 ;
  assign n22091 = x[2] & n22089 ;
  assign n30289 = ~n22091 ;
  assign n22092 = n22090 & n30289 ;
  assign n12749 = n3639 & n12695 ;
  assign n12671 = x[107] & n12633 ;
  assign n14377 = x[108] & n13533 ;
  assign n18803 = n12671 | n14377 ;
  assign n18804 = x[109] & n12631 ;
  assign n18805 = n18803 | n18804 ;
  assign n18806 = n12749 | n18805 ;
  assign n30290 = ~n18806 ;
  assign n18807 = x[11] & n30290 ;
  assign n18808 = n27892 & n18806 ;
  assign n18809 = n18807 | n18808 ;
  assign n15628 = n15625 & n15627 ;
  assign n15630 = n15625 | n15627 ;
  assign n30291 = ~n15628 ;
  assign n15631 = n30291 & n15630 ;
  assign n30292 = ~n16517 ;
  assign n16518 = n15631 & n30292 ;
  assign n30293 = ~n15631 ;
  assign n16614 = n30293 & n16517 ;
  assign n16615 = n16518 | n16614 ;
  assign n16623 = n16615 | n16622 ;
  assign n16624 = n16615 & n16622 ;
  assign n30294 = ~n16624 ;
  assign n17445 = n16623 & n30294 ;
  assign n30295 = ~n17173 ;
  assign n17446 = n30295 & n17445 ;
  assign n30296 = ~n17445 ;
  assign n17579 = n17173 & n30296 ;
  assign n17580 = n17446 | n17579 ;
  assign n17582 = n17576 & n17580 ;
  assign n18772 = n17582 | n18771 ;
  assign n16521 = n15628 | n16520 ;
  assign n15552 = n14630 | n15551 ;
  assign n2412 = n452 & n2410 ;
  assign n354 = x[92] & n330 ;
  assign n415 = x[93] & n390 ;
  assign n13710 = n354 | n415 ;
  assign n13711 = x[94] & n322 ;
  assign n13712 = n13710 | n13711 ;
  assign n13713 = n2412 | n13712 ;
  assign n30297 = ~n13713 ;
  assign n13714 = x[26] & n30297 ;
  assign n13715 = n28342 & n13713 ;
  assign n13716 = n13714 | n13715 ;
  assign n13429 = n13052 | n13428 ;
  assign n4665 = n2046 & n4632 ;
  assign n4515 = x[89] & n4514 ;
  assign n4577 = x[90] & n4572 ;
  assign n13033 = n4515 | n4577 ;
  assign n13034 = x[91] & n4504 ;
  assign n13035 = n13033 | n13034 ;
  assign n13036 = n4665 | n13035 ;
  assign n30298 = ~n13036 ;
  assign n13037 = x[29] & n30298 ;
  assign n13038 = n28483 & n13036 ;
  assign n13039 = n13037 | n13038 ;
  assign n12140 = n12137 & n12139 ;
  assign n30299 = ~n12205 ;
  assign n12208 = n12198 & n30299 ;
  assign n30300 = ~n12198 ;
  assign n12209 = n30300 & n12205 ;
  assign n12210 = n12208 | n12209 ;
  assign n12497 = n12210 & n12496 ;
  assign n12498 = n12207 | n12497 ;
  assign n12499 = n12196 & n12498 ;
  assign n12500 = n12195 | n12499 ;
  assign n12504 = n12500 & n12503 ;
  assign n12505 = n12140 | n12504 ;
  assign n1722 = n779 & n1720 ;
  assign n664 = x[86] & n663 ;
  assign n721 = x[87] & n720 ;
  assign n12121 = n664 | n721 ;
  assign n12122 = x[88] & n652 ;
  assign n12123 = n12121 | n12122 ;
  assign n12124 = n1722 | n12123 ;
  assign n30301 = ~n12124 ;
  assign n12125 = x[32] & n30301 ;
  assign n12126 = n28658 & n12124 ;
  assign n12127 = n12125 | n12126 ;
  assign n11411 = n11402 & n11409 ;
  assign n11686 = n11682 & n11684 ;
  assign n11687 = n11411 | n11686 ;
  assign n4053 = n1239 & n4041 ;
  assign n3933 = x[83] & n3910 ;
  assign n3998 = x[84] & n3975 ;
  assign n11389 = n3933 | n3998 ;
  assign n11390 = x[85] & n3906 ;
  assign n11391 = n11389 | n11390 ;
  assign n11392 = n4053 | n11391 ;
  assign n30302 = ~n11392 ;
  assign n11393 = x[35] & n30302 ;
  assign n11394 = n28822 & n11392 ;
  assign n11395 = n11393 | n11394 ;
  assign n10841 = n10838 & n10839 ;
  assign n11080 = n10841 | n11079 ;
  assign n3608 = n1003 & n3574 ;
  assign n3466 = x[80] & n3443 ;
  assign n3566 = x[81] & n3508 ;
  assign n10822 = n3466 | n3566 ;
  assign n10823 = x[82] & n3439 ;
  assign n10824 = n10822 | n10823 ;
  assign n10825 = n3608 | n10824 ;
  assign n30303 = ~n10825 ;
  assign n10826 = x[38] & n30303 ;
  assign n10827 = n28996 & n10825 ;
  assign n10828 = n10826 | n10827 ;
  assign n10126 = n30136 & n9620 ;
  assign n30304 = ~n9620 ;
  assign n10128 = n9618 & n30304 ;
  assign n10129 = n10126 | n10128 ;
  assign n10130 = n10125 & n10129 ;
  assign n10321 = n10130 | n10320 ;
  assign n3188 = n1741 & n3162 ;
  assign n3090 = x[77] & n3031 ;
  assign n3106 = x[78] & n3096 ;
  assign n10107 = n3090 | n3106 ;
  assign n10108 = x[79] & n3027 ;
  assign n10109 = n10107 | n10108 ;
  assign n10110 = n3188 | n10109 ;
  assign n30305 = ~n10110 ;
  assign n10111 = x[41] & n30305 ;
  assign n10112 = n29184 & n10110 ;
  assign n10113 = n10111 | n10112 ;
  assign n9478 = n9474 & n9476 ;
  assign n9622 = n9478 | n9621 ;
  assign n2754 = n2635 & n2750 ;
  assign n2522 = x[74] & n2492 ;
  assign n2587 = x[75] & n2557 ;
  assign n9458 = n2522 | n2587 ;
  assign n9459 = x[76] & n2488 ;
  assign n9460 = n9458 | n9459 ;
  assign n9461 = n2754 | n9460 ;
  assign n30306 = ~n9461 ;
  assign n9462 = x[44] & n30306 ;
  assign n9463 = n29400 & n9461 ;
  assign n9464 = n9462 | n9463 ;
  assign n9078 = n9075 | n9077 ;
  assign n3738 = n2321 & n3733 ;
  assign n2198 = x[71] & n2179 ;
  assign n2299 = x[72] & n2244 ;
  assign n8959 = n2198 | n2299 ;
  assign n8960 = x[73] & n2175 ;
  assign n8961 = n8959 | n8960 ;
  assign n8962 = n3738 | n8961 ;
  assign n30307 = ~n8962 ;
  assign n8963 = x[47] & n30307 ;
  assign n8964 = n29621 & n8962 ;
  assign n8965 = n8963 | n8964 ;
  assign n5984 = n2007 & n5976 ;
  assign n1892 = x[68] & n1866 ;
  assign n1952 = x[69] & n1931 ;
  assign n8365 = n1892 | n1952 ;
  assign n8366 = x[70] & n1862 ;
  assign n8367 = n8365 | n8366 ;
  assign n8368 = n5984 | n8367 ;
  assign n30308 = ~n8368 ;
  assign n8369 = x[50] & n30308 ;
  assign n8370 = n29865 & n8368 ;
  assign n8371 = n8369 | n8370 ;
  assign n27680 = x[53] & x[54] ;
  assign n1311 = x[53] | x[54] ;
  assign n30309 = ~n27680 ;
  assign n1312 = n30309 & n1311 ;
  assign n7398 = x[64] & n1312 ;
  assign n7933 = n7924 & n7931 ;
  assign n7934 = n7398 & n7933 ;
  assign n7935 = n7398 | n7933 ;
  assign n30310 = ~n7934 ;
  assign n7936 = n30310 & n7935 ;
  assign n6505 = n1690 & n6494 ;
  assign n1589 = x[65] & n1551 ;
  assign n1657 = x[66] & n1616 ;
  assign n7937 = n1589 | n1657 ;
  assign n7938 = x[67] & n1547 ;
  assign n7939 = n7937 | n7938 ;
  assign n7940 = n6505 | n7939 ;
  assign n30311 = ~n7940 ;
  assign n7941 = x[53] & n30311 ;
  assign n7942 = n30125 & n7940 ;
  assign n7943 = n7941 | n7942 ;
  assign n30312 = ~n7943 ;
  assign n7944 = n7936 & n30312 ;
  assign n30313 = ~n7936 ;
  assign n8372 = n30313 & n7943 ;
  assign n8373 = n7944 | n8372 ;
  assign n30314 = ~n8371 ;
  assign n8374 = n30314 & n8373 ;
  assign n30315 = ~n8373 ;
  assign n8438 = n8371 & n30315 ;
  assign n8439 = n8374 | n8438 ;
  assign n30316 = ~n8439 ;
  assign n8440 = n8437 & n30316 ;
  assign n8966 = n30226 & n8439 ;
  assign n8967 = n8440 | n8966 ;
  assign n30317 = ~n8967 ;
  assign n9079 = n8965 & n30317 ;
  assign n30318 = ~n8965 ;
  assign n9080 = n30318 & n8967 ;
  assign n9081 = n9079 | n9080 ;
  assign n9082 = n9078 & n9081 ;
  assign n9465 = n9078 | n9080 ;
  assign n9466 = n9079 | n9465 ;
  assign n30319 = ~n9082 ;
  assign n9467 = n30319 & n9466 ;
  assign n30320 = ~n9467 ;
  assign n9623 = n9464 & n30320 ;
  assign n30321 = ~n9464 ;
  assign n9624 = n30321 & n9467 ;
  assign n9625 = n9623 | n9624 ;
  assign n9626 = n9622 & n9625 ;
  assign n10114 = n9622 | n9624 ;
  assign n10115 = n9623 | n10114 ;
  assign n30322 = ~n9626 ;
  assign n10116 = n30322 & n10115 ;
  assign n10117 = n10113 | n10116 ;
  assign n10118 = n10113 & n10116 ;
  assign n30323 = ~n10118 ;
  assign n10322 = n10117 & n30323 ;
  assign n10323 = n10321 & n10322 ;
  assign n10829 = n10321 | n10322 ;
  assign n30324 = ~n10323 ;
  assign n10830 = n30324 & n10829 ;
  assign n30325 = ~n10828 ;
  assign n11081 = n30325 & n10830 ;
  assign n30326 = ~n10830 ;
  assign n11082 = n10828 & n30326 ;
  assign n11083 = n11081 | n11082 ;
  assign n11084 = n11080 & n11083 ;
  assign n11396 = n11080 | n11081 ;
  assign n11397 = n11082 | n11396 ;
  assign n30327 = ~n11084 ;
  assign n11398 = n30327 & n11397 ;
  assign n11399 = n11395 | n11398 ;
  assign n11400 = n11395 & n11398 ;
  assign n30328 = ~n11400 ;
  assign n11688 = n11399 & n30328 ;
  assign n11689 = n11687 & n11688 ;
  assign n12128 = n11687 | n11688 ;
  assign n30329 = ~n11689 ;
  assign n12129 = n30329 & n12128 ;
  assign n12130 = n12127 & n12129 ;
  assign n12506 = n12127 | n12129 ;
  assign n30330 = ~n12130 ;
  assign n12507 = n30330 & n12506 ;
  assign n12508 = n12505 & n12507 ;
  assign n13040 = n12505 | n12507 ;
  assign n30331 = ~n12508 ;
  assign n13041 = n30331 & n13040 ;
  assign n13042 = n13039 & n13041 ;
  assign n13430 = n13039 | n13041 ;
  assign n30332 = ~n13042 ;
  assign n13664 = n30332 & n13430 ;
  assign n30333 = ~n13429 ;
  assign n13666 = n30333 & n13664 ;
  assign n30334 = ~n13664 ;
  assign n13717 = n13429 & n30334 ;
  assign n13718 = n13666 | n13717 ;
  assign n30335 = ~n13716 ;
  assign n13719 = n30335 & n13718 ;
  assign n30336 = ~n13718 ;
  assign n14219 = n13716 & n30336 ;
  assign n14220 = n13719 | n14219 ;
  assign n14590 = n13832 & n13835 ;
  assign n14593 = n14195 & n14591 ;
  assign n14594 = n14590 | n14593 ;
  assign n14595 = n13814 | n13821 ;
  assign n14596 = n14594 & n14595 ;
  assign n14597 = n13823 | n14596 ;
  assign n14598 = n13746 | n13748 ;
  assign n30337 = ~n13749 ;
  assign n14599 = n30337 & n14598 ;
  assign n14600 = n14597 & n14599 ;
  assign n14601 = n13749 | n14600 ;
  assign n14602 = n13731 | n13738 ;
  assign n14603 = n14601 & n14602 ;
  assign n14604 = n14212 | n14603 ;
  assign n14606 = n14604 & n14605 ;
  assign n14608 = n13730 | n14606 ;
  assign n30338 = ~n14608 ;
  assign n14609 = n14220 & n30338 ;
  assign n30339 = ~n14220 ;
  assign n14610 = n30339 & n14608 ;
  assign n14611 = n14609 | n14610 ;
  assign n5327 = n2438 & n5302 ;
  assign n5264 = x[95] & n5240 ;
  assign n6275 = x[96] & n6179 ;
  assign n14612 = n5264 | n6275 ;
  assign n14613 = x[97] & n5238 ;
  assign n14614 = n14612 | n14613 ;
  assign n14615 = n5327 | n14614 ;
  assign n30340 = ~n14615 ;
  assign n14616 = x[23] & n30340 ;
  assign n14617 = n28221 & n14615 ;
  assign n14618 = n14616 | n14617 ;
  assign n30341 = ~n14618 ;
  assign n14619 = n14611 & n30341 ;
  assign n30342 = ~n14611 ;
  assign n15553 = n30342 & n14618 ;
  assign n15554 = n14619 | n15553 ;
  assign n15555 = n15552 | n15554 ;
  assign n15556 = n15552 & n15554 ;
  assign n30343 = ~n15556 ;
  assign n15609 = n15555 & n30343 ;
  assign n7218 = n2466 & n7162 ;
  assign n7134 = x[98] & n7100 ;
  assign n7690 = x[99] & n7647 ;
  assign n15610 = n7134 | n7690 ;
  assign n15611 = x[100] & n7098 ;
  assign n15612 = n15610 | n15611 ;
  assign n15613 = n7218 | n15612 ;
  assign n30344 = ~n15613 ;
  assign n15614 = x[20] & n30344 ;
  assign n15615 = n28114 & n15613 ;
  assign n15616 = n15614 | n15615 ;
  assign n15617 = n15609 | n15616 ;
  assign n15618 = n15609 & n15616 ;
  assign n30345 = ~n15618 ;
  assign n16522 = n15617 & n30345 ;
  assign n16523 = n16521 & n16522 ;
  assign n16601 = n16521 | n16522 ;
  assign n30346 = ~n16523 ;
  assign n16602 = n30346 & n16601 ;
  assign n8751 = n2626 & n8706 ;
  assign n8672 = x[101] & n8645 ;
  assign n9847 = x[102] & n9278 ;
  assign n16603 = n8672 | n9847 ;
  assign n16604 = x[103] & n8643 ;
  assign n16605 = n16603 | n16604 ;
  assign n16606 = n8751 | n16605 ;
  assign n30347 = ~n16606 ;
  assign n16607 = x[17] & n30347 ;
  assign n16608 = n28039 & n16606 ;
  assign n16609 = n16607 | n16608 ;
  assign n16611 = n16602 & n16609 ;
  assign n16612 = n16602 | n16609 ;
  assign n30348 = ~n16611 ;
  assign n16613 = n30348 & n16612 ;
  assign n17444 = n16622 & n16625 ;
  assign n17504 = n16642 | n17503 ;
  assign n17505 = n17445 & n17504 ;
  assign n17506 = n17444 | n17505 ;
  assign n30349 = ~n17506 ;
  assign n17507 = n16613 & n30349 ;
  assign n30350 = ~n16613 ;
  assign n17558 = n30350 & n17506 ;
  assign n17559 = n17507 | n17558 ;
  assign n10550 = n3223 & n10542 ;
  assign n10484 = x[104] & n10481 ;
  assign n11888 = x[105] & n11232 ;
  assign n17560 = n10484 | n11888 ;
  assign n17561 = x[106] & n10479 ;
  assign n17562 = n17560 | n17561 ;
  assign n17563 = n10550 | n17562 ;
  assign n30351 = ~n17563 ;
  assign n17564 = x[14] & n30351 ;
  assign n17565 = n27956 & n17563 ;
  assign n17566 = n17564 | n17565 ;
  assign n17567 = n17559 | n17566 ;
  assign n17568 = n17559 & n17566 ;
  assign n30352 = ~n17568 ;
  assign n18773 = n17567 & n30352 ;
  assign n18774 = n18772 & n18773 ;
  assign n18810 = n18772 | n18773 ;
  assign n30353 = ~n18774 ;
  assign n18811 = n30353 & n18810 ;
  assign n30354 = ~n18809 ;
  assign n18812 = n30354 & n18811 ;
  assign n30355 = ~n18811 ;
  assign n19549 = n18809 & n30355 ;
  assign n19550 = n18812 | n19549 ;
  assign n19551 = n19547 | n19550 ;
  assign n19552 = n19547 & n19550 ;
  assign n30356 = ~n19552 ;
  assign n20027 = n19551 & n30356 ;
  assign n15362 = n4442 & n15308 ;
  assign n15304 = x[110] & n15246 ;
  assign n17297 = x[111] & n16288 ;
  assign n20028 = n15304 | n17297 ;
  assign n20029 = x[112] & n15244 ;
  assign n20030 = n20028 | n20029 ;
  assign n20031 = n15362 | n20030 ;
  assign n30357 = ~n20031 ;
  assign n20032 = x[8] & n30357 ;
  assign n20033 = n27845 & n20031 ;
  assign n20034 = n20032 | n20033 ;
  assign n20035 = n20027 | n20034 ;
  assign n20036 = n20027 & n20034 ;
  assign n30358 = ~n20036 ;
  assign n20037 = n20035 & n30358 ;
  assign n20896 = n20123 | n20895 ;
  assign n20897 = n20037 | n20896 ;
  assign n20898 = n20037 & n20896 ;
  assign n30359 = ~n20898 ;
  assign n21068 = n20897 & n30359 ;
  assign n18411 = n4474 & n18392 ;
  assign n18385 = x[113] & n18329 ;
  assign n18518 = x[114] & n18514 ;
  assign n21069 = n18385 | n18518 ;
  assign n21070 = x[115] & n18327 ;
  assign n21071 = n21069 | n21070 ;
  assign n21072 = n18411 | n21071 ;
  assign n30360 = ~n21072 ;
  assign n21073 = x[5] & n30360 ;
  assign n21074 = n27813 & n21072 ;
  assign n21075 = n21073 | n21074 ;
  assign n21076 = n21068 | n21075 ;
  assign n21077 = n21068 & n21075 ;
  assign n30361 = ~n21077 ;
  assign n22016 = n21076 & n30361 ;
  assign n22017 = n22015 & n22016 ;
  assign n22093 = n22015 | n22016 ;
  assign n30362 = ~n22017 ;
  assign n22094 = n30362 & n22093 ;
  assign n22095 = n22092 & n22094 ;
  assign n23078 = n22092 | n22094 ;
  assign n30363 = ~n22095 ;
  assign n23079 = n30363 & n23078 ;
  assign n23080 = n23077 & n23079 ;
  assign n27702 = n23077 | n23079 ;
  assign n30364 = ~n23080 ;
  assign n183 = n30364 & n27702 ;
  assign n23081 = n22095 | n23080 ;
  assign n22018 = n21077 | n22017 ;
  assign n18440 = n4702 & n18392 ;
  assign n18356 = x[114] & n18329 ;
  assign n18571 = x[115] & n18514 ;
  assign n21057 = n18356 | n18571 ;
  assign n21058 = x[116] & n18327 ;
  assign n21059 = n21057 | n21058 ;
  assign n21060 = n18440 | n21059 ;
  assign n30365 = ~n21060 ;
  assign n21061 = x[5] & n30365 ;
  assign n21062 = n27813 & n21060 ;
  assign n21063 = n21061 | n21062 ;
  assign n20899 = n20036 | n20898 ;
  assign n15358 = n4087 & n15308 ;
  assign n15295 = x[111] & n15246 ;
  assign n17309 = x[112] & n16288 ;
  assign n20017 = n15295 | n17309 ;
  assign n20018 = x[113] & n15244 ;
  assign n20019 = n20017 | n20018 ;
  assign n20020 = n15358 | n20019 ;
  assign n20021 = x[8] | n20020 ;
  assign n20022 = x[8] & n20020 ;
  assign n30366 = ~n20022 ;
  assign n20023 = n20021 & n30366 ;
  assign n18813 = n18809 & n18811 ;
  assign n19553 = n18813 | n19552 ;
  assign n8737 = n3001 & n8706 ;
  assign n8679 = x[102] & n8645 ;
  assign n9848 = x[103] & n9278 ;
  assign n16588 = n8679 | n9848 ;
  assign n16589 = x[104] & n8643 ;
  assign n16590 = n16588 | n16589 ;
  assign n16591 = n8737 | n16590 ;
  assign n30367 = ~n16591 ;
  assign n16592 = x[17] & n30367 ;
  assign n16593 = n28039 & n16591 ;
  assign n16594 = n16592 | n16593 ;
  assign n3185 = n1270 & n3162 ;
  assign n3092 = x[78] & n3031 ;
  assign n3120 = x[79] & n3096 ;
  assign n10094 = n3092 | n3120 ;
  assign n10095 = x[80] & n3027 ;
  assign n10096 = n10094 | n10095 ;
  assign n10097 = n3185 | n10096 ;
  assign n30368 = ~n10097 ;
  assign n10098 = x[41] & n30368 ;
  assign n10099 = n29184 & n10097 ;
  assign n10100 = n10098 | n10099 ;
  assign n9627 = n9464 & n9467 ;
  assign n9628 = n9626 | n9627 ;
  assign n2640 = n1775 & n2635 ;
  assign n2506 = x[75] & n2492 ;
  assign n2586 = x[76] & n2557 ;
  assign n9448 = n2506 | n2586 ;
  assign n9449 = x[77] & n2488 ;
  assign n9450 = n9448 | n9449 ;
  assign n9451 = n2640 | n9450 ;
  assign n9452 = x[44] | n9451 ;
  assign n9453 = x[44] & n9451 ;
  assign n30369 = ~n9453 ;
  assign n9454 = n9452 & n30369 ;
  assign n8968 = n8965 & n8967 ;
  assign n9083 = n8968 | n9082 ;
  assign n2725 = n2321 & n2722 ;
  assign n2194 = x[72] & n2179 ;
  assign n2270 = x[73] & n2244 ;
  assign n8948 = n2194 | n2270 ;
  assign n8949 = x[74] & n2175 ;
  assign n8950 = n8948 | n8949 ;
  assign n8951 = n2725 | n8950 ;
  assign n30370 = ~n8951 ;
  assign n8952 = x[47] & n30370 ;
  assign n8953 = n29621 & n8951 ;
  assign n8954 = n8952 | n8953 ;
  assign n8375 = n8371 & n8373 ;
  assign n8441 = n8437 & n8439 ;
  assign n8442 = n8375 | n8441 ;
  assign n4793 = n2007 & n4790 ;
  assign n1893 = x[69] & n1866 ;
  assign n1954 = x[70] & n1931 ;
  assign n8354 = n1893 | n1954 ;
  assign n8355 = x[71] & n1862 ;
  assign n8356 = n8354 | n8355 ;
  assign n8357 = n4793 | n8356 ;
  assign n30371 = ~n8357 ;
  assign n8358 = x[50] & n30371 ;
  assign n8359 = n29865 & n8357 ;
  assign n8360 = n8358 | n8359 ;
  assign n7945 = n7936 & n7943 ;
  assign n7946 = n7934 | n7945 ;
  assign n6421 = n1690 & n6408 ;
  assign n1574 = x[66] & n1551 ;
  assign n1634 = x[67] & n1616 ;
  assign n7903 = n1574 | n1634 ;
  assign n7904 = x[68] & n1547 ;
  assign n7905 = n7903 | n7904 ;
  assign n7906 = n6421 | n7905 ;
  assign n30372 = ~n7906 ;
  assign n7907 = x[53] & n30372 ;
  assign n7908 = n30125 & n7906 ;
  assign n7909 = n7907 | n7908 ;
  assign n30373 = ~n7398 ;
  assign n7399 = x[56] & n30373 ;
  assign n27682 = x[55] & x[56] ;
  assign n1313 = x[55] | x[56] ;
  assign n30374 = ~n27682 ;
  assign n1314 = n30374 & n1313 ;
  assign n1457 = n1312 & n1314 ;
  assign n6448 = n1457 & n6437 ;
  assign n30375 = ~n1314 ;
  assign n1315 = n1312 & n30375 ;
  assign n7400 = x[65] & n1315 ;
  assign n27683 = x[54] & x[55] ;
  assign n1316 = x[54] | x[55] ;
  assign n30376 = ~n27683 ;
  assign n1317 = n30376 & n1316 ;
  assign n30377 = ~n1312 ;
  assign n1384 = n30377 & n1317 ;
  assign n7401 = x[64] & n1384 ;
  assign n7402 = n7400 | n7401 ;
  assign n7403 = n6448 | n7402 ;
  assign n30378 = ~n7403 ;
  assign n7404 = x[56] & n30378 ;
  assign n30379 = ~x[56] ;
  assign n7405 = n30379 & n7403 ;
  assign n7406 = n7404 | n7405 ;
  assign n30380 = ~n7406 ;
  assign n7407 = n7399 & n30380 ;
  assign n30381 = ~n7399 ;
  assign n7910 = n30381 & n7406 ;
  assign n7911 = n7407 | n7910 ;
  assign n30382 = ~n7909 ;
  assign n7912 = n30382 & n7911 ;
  assign n30383 = ~n7911 ;
  assign n7947 = n7909 & n30383 ;
  assign n7948 = n7912 | n7947 ;
  assign n30384 = ~n7946 ;
  assign n7949 = n30384 & n7948 ;
  assign n30385 = ~n7948 ;
  assign n8361 = n7946 & n30385 ;
  assign n8362 = n7949 | n8361 ;
  assign n30386 = ~n8360 ;
  assign n8363 = n30386 & n8362 ;
  assign n30387 = ~n8362 ;
  assign n8443 = n8360 & n30387 ;
  assign n8444 = n8363 | n8443 ;
  assign n30388 = ~n8442 ;
  assign n8445 = n30388 & n8444 ;
  assign n30389 = ~n8444 ;
  assign n8955 = n8442 & n30389 ;
  assign n8956 = n8445 | n8955 ;
  assign n30390 = ~n8954 ;
  assign n8957 = n30390 & n8956 ;
  assign n30391 = ~n8956 ;
  assign n9084 = n8954 & n30391 ;
  assign n9085 = n8957 | n9084 ;
  assign n30392 = ~n9083 ;
  assign n9086 = n30392 & n9085 ;
  assign n30393 = ~n9085 ;
  assign n9455 = n9083 & n30393 ;
  assign n9456 = n9086 | n9455 ;
  assign n9457 = n9454 & n9456 ;
  assign n9629 = n9454 | n9456 ;
  assign n30394 = ~n9457 ;
  assign n9630 = n30394 & n9629 ;
  assign n9631 = n9628 & n9630 ;
  assign n10101 = n9628 | n9630 ;
  assign n30395 = ~n9631 ;
  assign n10102 = n30395 & n10101 ;
  assign n30396 = ~n10100 ;
  assign n10104 = n30396 & n10102 ;
  assign n30397 = ~n10102 ;
  assign n10105 = n10100 & n30397 ;
  assign n10106 = n10104 | n10105 ;
  assign n10324 = n10118 | n10323 ;
  assign n10325 = n10106 | n10324 ;
  assign n10326 = n10106 & n10324 ;
  assign n30398 = ~n10326 ;
  assign n10813 = n10325 & n30398 ;
  assign n3582 = n1057 & n3574 ;
  assign n3467 = x[81] & n3443 ;
  assign n3557 = x[82] & n3508 ;
  assign n10814 = n3467 | n3557 ;
  assign n10815 = x[83] & n3439 ;
  assign n10816 = n10814 | n10815 ;
  assign n10817 = n3582 | n10816 ;
  assign n30399 = ~n10817 ;
  assign n10818 = x[38] & n30399 ;
  assign n10819 = n28996 & n10817 ;
  assign n10820 = n10818 | n10819 ;
  assign n11086 = n10813 | n10820 ;
  assign n10821 = n10813 & n10820 ;
  assign n10831 = n10828 & n10830 ;
  assign n11085 = n10831 | n11084 ;
  assign n11087 = n11085 & n11086 ;
  assign n11088 = n10821 | n11087 ;
  assign n30400 = ~n11088 ;
  assign n11089 = n11086 & n30400 ;
  assign n30401 = ~n10821 ;
  assign n11376 = n30401 & n11086 ;
  assign n30402 = ~n11376 ;
  assign n11377 = n11085 & n30402 ;
  assign n11378 = n11089 | n11377 ;
  assign n4043 = n1213 & n4041 ;
  assign n3934 = x[84] & n3910 ;
  assign n4000 = x[85] & n3975 ;
  assign n11379 = n3934 | n4000 ;
  assign n11380 = x[86] & n3906 ;
  assign n11381 = n11379 | n11380 ;
  assign n11382 = n4043 | n11381 ;
  assign n30403 = ~n11382 ;
  assign n11383 = x[35] & n30403 ;
  assign n11384 = n28822 & n11382 ;
  assign n11385 = n11383 | n11384 ;
  assign n11386 = n11378 | n11385 ;
  assign n11387 = n11378 & n11385 ;
  assign n30404 = ~n11387 ;
  assign n11388 = n11386 & n30404 ;
  assign n11690 = n11400 | n11689 ;
  assign n11691 = n11388 | n11690 ;
  assign n11692 = n11388 & n11690 ;
  assign n30405 = ~n11692 ;
  assign n12108 = n11691 & n30405 ;
  assign n1456 = n779 & n1453 ;
  assign n666 = x[87] & n663 ;
  assign n722 = x[88] & n720 ;
  assign n12109 = n666 | n722 ;
  assign n12110 = x[89] & n652 ;
  assign n12111 = n12109 | n12110 ;
  assign n12112 = n1456 | n12111 ;
  assign n30406 = ~n12112 ;
  assign n12113 = x[32] & n30406 ;
  assign n12114 = n28658 & n12112 ;
  assign n12115 = n12113 | n12114 ;
  assign n30407 = ~n12115 ;
  assign n12118 = n12108 & n30407 ;
  assign n30408 = ~n12108 ;
  assign n12119 = n30408 & n12115 ;
  assign n12120 = n12118 | n12119 ;
  assign n12509 = n12130 | n12508 ;
  assign n12510 = n12120 | n12509 ;
  assign n12511 = n12120 & n12509 ;
  assign n30409 = ~n12511 ;
  assign n13018 = n12510 & n30409 ;
  assign n4657 = n1841 & n4632 ;
  assign n4544 = x[90] & n4514 ;
  assign n4582 = x[91] & n4572 ;
  assign n13019 = n4544 | n4582 ;
  assign n13020 = x[92] & n4504 ;
  assign n13021 = n13019 | n13020 ;
  assign n13022 = n4657 | n13021 ;
  assign n30410 = ~n13022 ;
  assign n13023 = x[29] & n30410 ;
  assign n13024 = n28483 & n13022 ;
  assign n13025 = n13023 | n13024 ;
  assign n30411 = ~n13025 ;
  assign n13026 = n13018 & n30411 ;
  assign n30412 = ~n13018 ;
  assign n13655 = n30412 & n13025 ;
  assign n13656 = n13026 | n13655 ;
  assign n13657 = n13061 & n13419 ;
  assign n13062 = n13054 | n13061 ;
  assign n30413 = ~n13063 ;
  assign n13659 = n13062 & n30413 ;
  assign n13660 = n13418 & n13659 ;
  assign n13661 = n13657 | n13660 ;
  assign n13662 = n13426 & n13661 ;
  assign n13663 = n13052 | n13662 ;
  assign n13665 = n13663 & n13664 ;
  assign n13667 = n13042 | n13665 ;
  assign n13668 = n13656 | n13667 ;
  assign n13669 = n13656 & n13667 ;
  assign n30414 = ~n13669 ;
  assign n13698 = n13668 & n30414 ;
  assign n2153 = n452 & n2152 ;
  assign n357 = x[93] & n330 ;
  assign n414 = x[94] & n390 ;
  assign n13699 = n357 | n414 ;
  assign n13700 = x[95] & n322 ;
  assign n13701 = n13699 | n13700 ;
  assign n13702 = n2153 | n13701 ;
  assign n30415 = ~n13702 ;
  assign n13703 = x[26] & n30415 ;
  assign n13704 = n28342 & n13702 ;
  assign n13705 = n13703 | n13704 ;
  assign n30416 = ~n13705 ;
  assign n13706 = n13698 & n30416 ;
  assign n30417 = ~n13698 ;
  assign n13708 = n30417 & n13705 ;
  assign n13709 = n13706 | n13708 ;
  assign n13720 = n13716 & n13718 ;
  assign n14217 = n14215 & n14216 ;
  assign n14218 = n13730 | n14217 ;
  assign n14221 = n14218 & n14220 ;
  assign n14222 = n13720 | n14221 ;
  assign n14223 = n13709 | n14222 ;
  assign n14224 = n13709 & n14222 ;
  assign n30418 = ~n14224 ;
  assign n14577 = n14223 & n30418 ;
  assign n5328 = n2841 & n5302 ;
  assign n5299 = x[96] & n5240 ;
  assign n6269 = x[97] & n6179 ;
  assign n14578 = n5299 | n6269 ;
  assign n14579 = x[98] & n5238 ;
  assign n14580 = n14578 | n14579 ;
  assign n14581 = n5328 | n14580 ;
  assign n30419 = ~n14581 ;
  assign n14582 = x[23] & n30419 ;
  assign n14583 = n28221 & n14581 ;
  assign n14584 = n14582 | n14583 ;
  assign n30420 = ~n14584 ;
  assign n14587 = n14577 & n30420 ;
  assign n30421 = ~n14577 ;
  assign n14588 = n30421 & n14584 ;
  assign n14589 = n14587 | n14588 ;
  assign n14620 = n14611 & n14618 ;
  assign n15145 = n14652 & n15144 ;
  assign n15146 = n14653 | n15145 ;
  assign n15147 = n14643 & n15146 ;
  assign n15148 = n14641 | n15147 ;
  assign n15150 = n15148 & n15149 ;
  assign n15151 = n14630 | n15150 ;
  assign n15152 = n14611 | n14618 ;
  assign n30422 = ~n14620 ;
  assign n15153 = n30422 & n15152 ;
  assign n15154 = n15151 & n15153 ;
  assign n15155 = n14620 | n15154 ;
  assign n15156 = n14589 | n15155 ;
  assign n15157 = n14589 & n15155 ;
  assign n30423 = ~n15157 ;
  assign n15594 = n15156 & n30423 ;
  assign n7203 = n2977 & n7162 ;
  assign n7139 = x[99] & n7100 ;
  assign n7708 = x[100] & n7647 ;
  assign n15595 = n7139 | n7708 ;
  assign n15596 = x[101] & n7098 ;
  assign n15597 = n15595 | n15596 ;
  assign n15598 = n7203 | n15597 ;
  assign n30424 = ~n15598 ;
  assign n15599 = x[20] & n30424 ;
  assign n15600 = n28114 & n15598 ;
  assign n15601 = n15599 | n15600 ;
  assign n30425 = ~n15601 ;
  assign n15602 = n15594 & n30425 ;
  assign n30426 = ~n15594 ;
  assign n16393 = n30426 & n15601 ;
  assign n16394 = n15602 | n16393 ;
  assign n16524 = n15618 | n16523 ;
  assign n16526 = n16394 | n16524 ;
  assign n16527 = n16394 & n16524 ;
  assign n30427 = ~n16527 ;
  assign n16597 = n16526 & n30427 ;
  assign n30428 = ~n16594 ;
  assign n16598 = n30428 & n16597 ;
  assign n30429 = ~n16597 ;
  assign n16599 = n16594 & n30429 ;
  assign n16600 = n16598 | n16599 ;
  assign n17176 = n16624 | n17175 ;
  assign n17177 = n16613 & n17176 ;
  assign n17178 = n16611 | n17177 ;
  assign n17179 = n16600 | n17178 ;
  assign n17180 = n16600 & n17178 ;
  assign n30430 = ~n17180 ;
  assign n17549 = n17179 & n30430 ;
  assign n10574 = n3199 & n10542 ;
  assign n10485 = x[105] & n10481 ;
  assign n11877 = x[106] & n11232 ;
  assign n17550 = n10485 | n11877 ;
  assign n17551 = x[107] & n10479 ;
  assign n17552 = n17550 | n17551 ;
  assign n17553 = n10574 | n17552 ;
  assign n30431 = ~n17553 ;
  assign n17554 = x[14] & n30431 ;
  assign n17555 = n27956 & n17553 ;
  assign n17556 = n17554 | n17555 ;
  assign n18254 = n17549 | n17556 ;
  assign n17557 = n17549 & n17556 ;
  assign n17578 = n17569 & n17576 ;
  assign n17581 = n17576 | n17580 ;
  assign n30432 = ~n17582 ;
  assign n17583 = n17581 & n30432 ;
  assign n18247 = n17594 | n18246 ;
  assign n18248 = n17583 & n18247 ;
  assign n18249 = n17578 | n18248 ;
  assign n30433 = ~n16609 ;
  assign n16610 = n16602 & n30433 ;
  assign n30434 = ~n16602 ;
  assign n17442 = n30434 & n16609 ;
  assign n17443 = n16610 | n17442 ;
  assign n17508 = n17443 | n17506 ;
  assign n17509 = n17443 & n17506 ;
  assign n30435 = ~n17509 ;
  assign n18250 = n17508 & n30435 ;
  assign n18251 = n17566 | n18250 ;
  assign n18252 = n18249 & n18251 ;
  assign n18253 = n17568 | n18252 ;
  assign n18255 = n18253 & n18254 ;
  assign n18256 = n17557 | n18255 ;
  assign n30436 = ~n18256 ;
  assign n18257 = n18254 & n30436 ;
  assign n18684 = n17566 & n18250 ;
  assign n18775 = n18684 | n18774 ;
  assign n30437 = ~n17557 ;
  assign n18791 = n30437 & n18254 ;
  assign n30438 = ~n18791 ;
  assign n18792 = n18775 & n30438 ;
  assign n18793 = n18257 | n18792 ;
  assign n12748 = n3615 & n12695 ;
  assign n12678 = x[108] & n12633 ;
  assign n14394 = x[109] & n13533 ;
  assign n18794 = n12678 | n14394 ;
  assign n18795 = x[110] & n12631 ;
  assign n18796 = n18794 | n18795 ;
  assign n18797 = n12748 | n18796 ;
  assign n30439 = ~n18797 ;
  assign n18798 = x[11] & n30439 ;
  assign n18799 = n27892 & n18797 ;
  assign n18800 = n18798 | n18799 ;
  assign n18801 = n18793 | n18800 ;
  assign n18802 = n18793 & n18800 ;
  assign n30440 = ~n18802 ;
  assign n19554 = n18801 & n30440 ;
  assign n19555 = n19553 & n19554 ;
  assign n20024 = n19553 | n19554 ;
  assign n30441 = ~n19555 ;
  assign n20025 = n30441 & n20024 ;
  assign n20026 = n20023 & n20025 ;
  assign n20900 = n20023 | n20025 ;
  assign n30442 = ~n20026 ;
  assign n20901 = n30442 & n20900 ;
  assign n20902 = n20899 & n20901 ;
  assign n21064 = n20899 | n20901 ;
  assign n30443 = ~n20902 ;
  assign n21065 = n30443 & n21064 ;
  assign n30444 = ~n21063 ;
  assign n21066 = n30444 & n21065 ;
  assign n30445 = ~n21065 ;
  assign n22019 = n21063 & n30445 ;
  assign n22020 = n21066 | n22019 ;
  assign n22021 = n22018 | n22020 ;
  assign n22022 = n22018 & n22020 ;
  assign n30446 = ~n22022 ;
  assign n22076 = n22021 & n30446 ;
  assign n618 = n616 & n617 ;
  assign n619 = n24007 | n618 ;
  assign n27542 = x[118] & x[119] ;
  assign n620 = x[118] | x[119] ;
  assign n30447 = ~n27542 ;
  assign n5044 = n30447 & n620 ;
  assign n5045 = n619 | n5044 ;
  assign n5046 = n619 & n5044 ;
  assign n30448 = ~n5046 ;
  assign n5047 = n5045 & n30448 ;
  assign n19677 = n5047 & n19656 ;
  assign n19751 = x[117] & n19723 ;
  assign n19875 = x[118] & n19829 ;
  assign n22077 = n19751 | n19875 ;
  assign n22078 = x[119] & n19655 ;
  assign n22079 = n22077 | n22078 ;
  assign n22080 = n19677 | n22079 ;
  assign n30449 = ~n22080 ;
  assign n22081 = x[2] & n30449 ;
  assign n22082 = n27790 & n22080 ;
  assign n22083 = n22081 | n22082 ;
  assign n22084 = n22076 | n22083 ;
  assign n22085 = n22076 & n22083 ;
  assign n30450 = ~n22085 ;
  assign n23082 = n22084 & n30450 ;
  assign n23083 = n23081 | n23082 ;
  assign n23084 = n23081 & n23082 ;
  assign n30451 = ~n23084 ;
  assign n184 = n23083 & n30451 ;
  assign n621 = n619 & n620 ;
  assign n622 = n27542 | n621 ;
  assign n23813 = x[119] & x[120] ;
  assign n623 = x[119] | x[120] ;
  assign n30452 = ~n23813 ;
  assign n4675 = n30452 & n623 ;
  assign n4676 = n622 & n4675 ;
  assign n4677 = n622 | n4675 ;
  assign n30453 = ~n4676 ;
  assign n4678 = n30453 & n4677 ;
  assign n19681 = n4678 & n19656 ;
  assign n19766 = x[118] & n19723 ;
  assign n19859 = x[119] & n19829 ;
  assign n22064 = n19766 | n19859 ;
  assign n22065 = x[120] & n19655 ;
  assign n22066 = n22064 | n22065 ;
  assign n22067 = n19681 | n22066 ;
  assign n22068 = x[2] | n22067 ;
  assign n22069 = x[2] & n22067 ;
  assign n30454 = ~n22069 ;
  assign n22070 = n22068 & n30454 ;
  assign n21067 = n21063 & n21065 ;
  assign n22023 = n21067 | n22022 ;
  assign n20903 = n20026 | n20902 ;
  assign n15366 = n4276 & n15308 ;
  assign n15290 = x[112] & n15246 ;
  assign n17304 = x[113] & n16288 ;
  assign n20007 = n15290 | n17304 ;
  assign n20008 = x[114] & n15244 ;
  assign n20009 = n20007 | n20008 ;
  assign n20010 = n15366 | n20009 ;
  assign n30455 = ~n20010 ;
  assign n20011 = x[8] & n30455 ;
  assign n20012 = n27845 & n20010 ;
  assign n20013 = n20011 | n20012 ;
  assign n19556 = n18802 | n19555 ;
  assign n18776 = n18254 & n18775 ;
  assign n18777 = n17557 | n18776 ;
  assign n8748 = n3409 & n8706 ;
  assign n8700 = x[103] & n8645 ;
  assign n9849 = x[104] & n9278 ;
  assign n16572 = n8700 | n9849 ;
  assign n16573 = x[105] & n8643 ;
  assign n16574 = n16572 | n16573 ;
  assign n16575 = n8748 | n16574 ;
  assign n30456 = ~n16575 ;
  assign n16576 = x[17] & n30456 ;
  assign n16577 = n28039 & n16575 ;
  assign n16578 = n16576 | n16577 ;
  assign n15603 = n15594 & n15601 ;
  assign n14585 = n14577 | n14584 ;
  assign n14586 = n14577 & n14584 ;
  assign n30457 = ~n14586 ;
  assign n15516 = n14585 & n30457 ;
  assign n30458 = ~n15155 ;
  assign n15517 = n30458 & n15516 ;
  assign n30459 = ~n15516 ;
  assign n15604 = n15155 & n30459 ;
  assign n15605 = n15517 | n15604 ;
  assign n15606 = n15601 | n15605 ;
  assign n15607 = n15601 & n15605 ;
  assign n30460 = ~n15607 ;
  assign n15608 = n15606 & n30460 ;
  assign n16212 = n15642 | n16211 ;
  assign n16213 = n15631 & n16212 ;
  assign n16214 = n15628 | n16213 ;
  assign n16215 = n15617 & n16214 ;
  assign n16216 = n15618 | n16215 ;
  assign n16217 = n15608 & n16216 ;
  assign n16218 = n15603 | n16217 ;
  assign n5342 = n2313 & n5302 ;
  assign n5275 = x[97] & n5240 ;
  assign n6235 = x[98] & n6179 ;
  assign n14564 = n5275 | n6235 ;
  assign n14565 = x[99] & n5238 ;
  assign n14566 = n14564 | n14565 ;
  assign n14567 = n5342 | n14566 ;
  assign n30461 = ~n14567 ;
  assign n14568 = x[23] & n30461 ;
  assign n14569 = n28221 & n14567 ;
  assign n14570 = n14568 | n14569 ;
  assign n13707 = n13698 & n13705 ;
  assign n14225 = n13707 | n14224 ;
  assign n2001 = n452 & n2000 ;
  assign n388 = x[94] & n330 ;
  assign n391 = x[95] & n390 ;
  assign n13687 = n388 | n391 ;
  assign n13688 = x[96] & n322 ;
  assign n13689 = n13687 | n13688 ;
  assign n13690 = n2001 | n13689 ;
  assign n30462 = ~n13690 ;
  assign n13691 = x[26] & n30462 ;
  assign n13692 = n28342 & n13690 ;
  assign n13693 = n13691 | n13692 ;
  assign n12116 = n12108 | n12115 ;
  assign n12117 = n12108 & n12115 ;
  assign n30463 = ~n12117 ;
  assign n12852 = n12116 & n30463 ;
  assign n30464 = ~n12509 ;
  assign n12853 = n30464 & n12852 ;
  assign n30465 = ~n12852 ;
  assign n13028 = n12509 & n30465 ;
  assign n13029 = n12853 | n13028 ;
  assign n13031 = n13025 & n13029 ;
  assign n13670 = n13031 | n13669 ;
  assign n12512 = n12117 | n12511 ;
  assign n11693 = n11387 | n11692 ;
  assign n10103 = n10100 & n10102 ;
  assign n10327 = n10103 | n10326 ;
  assign n3169 = n1029 & n3162 ;
  assign n3056 = x[79] & n3031 ;
  assign n3121 = x[80] & n3096 ;
  assign n10085 = n3056 | n3121 ;
  assign n10086 = x[81] & n3027 ;
  assign n10087 = n10085 | n10086 ;
  assign n10088 = n3169 | n10087 ;
  assign n30466 = ~n10088 ;
  assign n10089 = x[41] & n30466 ;
  assign n10090 = n29184 & n10088 ;
  assign n10091 = n10089 | n10090 ;
  assign n9632 = n9457 | n9631 ;
  assign n2638 = n2084 & n2635 ;
  assign n2507 = x[76] & n2492 ;
  assign n2584 = x[77] & n2557 ;
  assign n9437 = n2507 | n2584 ;
  assign n9438 = x[78] & n2488 ;
  assign n9439 = n9437 | n9438 ;
  assign n9440 = n2638 | n9439 ;
  assign n30467 = ~n9440 ;
  assign n9441 = x[44] & n30467 ;
  assign n9442 = n29400 & n9440 ;
  assign n9443 = n9441 | n9442 ;
  assign n8958 = n8954 & n8956 ;
  assign n9087 = n9083 & n9085 ;
  assign n9088 = n8958 | n9087 ;
  assign n3296 = n2321 & n3289 ;
  assign n2237 = x[73] & n2179 ;
  assign n2272 = x[74] & n2244 ;
  assign n8937 = n2237 | n2272 ;
  assign n8938 = x[75] & n2175 ;
  assign n8939 = n8937 | n8938 ;
  assign n8940 = n3296 | n8939 ;
  assign n30468 = ~n8940 ;
  assign n8941 = x[47] & n30468 ;
  assign n8942 = n29621 & n8940 ;
  assign n8943 = n8941 | n8942 ;
  assign n8364 = n8360 & n8362 ;
  assign n8446 = n8442 & n8444 ;
  assign n8447 = n8364 | n8446 ;
  assign n7408 = n7399 & n7406 ;
  assign n6476 = n1457 & n6466 ;
  assign n1318 = n30377 & n1314 ;
  assign n30469 = ~n1317 ;
  assign n1319 = n30469 & n1318 ;
  assign n1345 = x[64] & n1319 ;
  assign n1436 = x[65] & n1384 ;
  assign n7409 = n1345 | n1436 ;
  assign n7410 = x[66] & n1315 ;
  assign n7411 = n7409 | n7410 ;
  assign n7412 = n6476 | n7411 ;
  assign n30470 = ~n7412 ;
  assign n7413 = x[56] & n30470 ;
  assign n7414 = n30379 & n7412 ;
  assign n7415 = n7413 | n7414 ;
  assign n30471 = ~n7415 ;
  assign n7416 = n7408 & n30471 ;
  assign n30472 = ~n7408 ;
  assign n7893 = n30472 & n7415 ;
  assign n7894 = n7416 | n7893 ;
  assign n6386 = n1690 & n6379 ;
  assign n1609 = x[67] & n1551 ;
  assign n1636 = x[68] & n1616 ;
  assign n7895 = n1609 | n1636 ;
  assign n7896 = x[69] & n1547 ;
  assign n7897 = n7895 | n7896 ;
  assign n7898 = n6386 | n7897 ;
  assign n30473 = ~n7898 ;
  assign n7899 = x[53] & n30473 ;
  assign n7900 = n30125 & n7898 ;
  assign n7901 = n7899 | n7900 ;
  assign n7952 = n7894 | n7901 ;
  assign n7902 = n7894 & n7901 ;
  assign n7913 = n7909 & n7911 ;
  assign n7950 = n7946 & n7948 ;
  assign n7951 = n7913 | n7950 ;
  assign n7954 = n7951 & n7952 ;
  assign n7955 = n7902 | n7954 ;
  assign n30474 = ~n7955 ;
  assign n7956 = n7952 & n30474 ;
  assign n30475 = ~n7902 ;
  assign n7953 = n30475 & n7952 ;
  assign n30476 = ~n7953 ;
  assign n8344 = n7951 & n30476 ;
  assign n8345 = n7956 | n8344 ;
  assign n3707 = n2007 & n3701 ;
  assign n1894 = x[70] & n1866 ;
  assign n1955 = x[71] & n1931 ;
  assign n8346 = n1894 | n1955 ;
  assign n8347 = x[72] & n1862 ;
  assign n8348 = n8346 | n8347 ;
  assign n8349 = n3707 | n8348 ;
  assign n30477 = ~n8349 ;
  assign n8350 = x[50] & n30477 ;
  assign n8351 = n29865 & n8349 ;
  assign n8352 = n8350 | n8351 ;
  assign n8353 = n8345 | n8352 ;
  assign n8448 = n8345 & n8352 ;
  assign n30478 = ~n8448 ;
  assign n8449 = n8353 & n30478 ;
  assign n30479 = ~n8447 ;
  assign n8450 = n30479 & n8449 ;
  assign n30480 = ~n8449 ;
  assign n8944 = n8447 & n30480 ;
  assign n8945 = n8450 | n8944 ;
  assign n30481 = ~n8943 ;
  assign n8946 = n30481 & n8945 ;
  assign n30482 = ~n8945 ;
  assign n9089 = n8943 & n30482 ;
  assign n9090 = n8946 | n9089 ;
  assign n9091 = n9088 & n9090 ;
  assign n9444 = n9088 | n9090 ;
  assign n30483 = ~n9091 ;
  assign n9445 = n30483 & n9444 ;
  assign n30484 = ~n9443 ;
  assign n9446 = n30484 & n9445 ;
  assign n30485 = ~n9445 ;
  assign n9633 = n9443 & n30485 ;
  assign n9634 = n9446 | n9633 ;
  assign n9635 = n9632 | n9634 ;
  assign n9636 = n9632 & n9634 ;
  assign n30486 = ~n9636 ;
  assign n10092 = n9635 & n30486 ;
  assign n30487 = ~n10091 ;
  assign n10328 = n30487 & n10092 ;
  assign n30488 = ~n10092 ;
  assign n10763 = n10091 & n30488 ;
  assign n10764 = n10328 | n10763 ;
  assign n30489 = ~n10764 ;
  assign n10765 = n10327 & n30489 ;
  assign n30490 = ~n10327 ;
  assign n10802 = n30490 & n10764 ;
  assign n10803 = n10765 | n10802 ;
  assign n3585 = n1293 & n3574 ;
  assign n3468 = x[82] & n3443 ;
  assign n3521 = x[83] & n3508 ;
  assign n10804 = n3468 | n3521 ;
  assign n10805 = x[84] & n3439 ;
  assign n10806 = n10804 | n10805 ;
  assign n10807 = n3585 | n10806 ;
  assign n30491 = ~n10807 ;
  assign n10808 = x[38] & n30491 ;
  assign n10809 = n28996 & n10807 ;
  assign n10810 = n10808 | n10809 ;
  assign n30492 = ~n10810 ;
  assign n10811 = n10803 & n30492 ;
  assign n30493 = ~n10803 ;
  assign n11090 = n30493 & n10810 ;
  assign n11091 = n10811 | n11090 ;
  assign n11092 = n11088 | n11091 ;
  assign n11093 = n11088 & n11091 ;
  assign n30494 = ~n11093 ;
  assign n11367 = n11092 & n30494 ;
  assign n4046 = n1522 & n4041 ;
  assign n3966 = x[85] & n3910 ;
  assign n4003 = x[86] & n3975 ;
  assign n11368 = n3966 | n4003 ;
  assign n11369 = x[87] & n3906 ;
  assign n11370 = n11368 | n11369 ;
  assign n11371 = n4046 | n11370 ;
  assign n30495 = ~n11371 ;
  assign n11372 = x[35] & n30495 ;
  assign n11373 = n28822 & n11371 ;
  assign n11374 = n11372 | n11373 ;
  assign n11375 = n11367 & n11374 ;
  assign n11694 = n11367 | n11374 ;
  assign n30496 = ~n11375 ;
  assign n11695 = n30496 & n11694 ;
  assign n11696 = n11693 & n11695 ;
  assign n12098 = n11693 | n11695 ;
  assign n30497 = ~n11696 ;
  assign n12099 = n30497 & n12098 ;
  assign n1483 = n779 & n1482 ;
  assign n689 = x[88] & n663 ;
  assign n723 = x[89] & n720 ;
  assign n12100 = n689 | n723 ;
  assign n12101 = x[90] & n652 ;
  assign n12102 = n12100 | n12101 ;
  assign n12103 = n1483 | n12102 ;
  assign n30498 = ~n12103 ;
  assign n12104 = x[32] & n30498 ;
  assign n12105 = n28658 & n12103 ;
  assign n12106 = n12104 | n12105 ;
  assign n12107 = n12099 & n12106 ;
  assign n12513 = n12099 | n12106 ;
  assign n30499 = ~n12107 ;
  assign n13005 = n30499 & n12513 ;
  assign n30500 = ~n13005 ;
  assign n13006 = n12512 & n30500 ;
  assign n12907 = n12137 | n12139 ;
  assign n30501 = ~n12140 ;
  assign n12908 = n30501 & n12907 ;
  assign n12909 = n12905 & n12908 ;
  assign n12910 = n12140 | n12909 ;
  assign n12911 = n12506 & n12910 ;
  assign n12912 = n12130 | n12911 ;
  assign n12913 = n12852 & n12912 ;
  assign n12914 = n12117 | n12913 ;
  assign n12915 = n12513 & n12914 ;
  assign n12916 = n12107 | n12915 ;
  assign n30502 = ~n12916 ;
  assign n13007 = n12513 & n30502 ;
  assign n13008 = n13006 | n13007 ;
  assign n4672 = n1685 & n4632 ;
  assign n4547 = x[91] & n4514 ;
  assign n4579 = x[92] & n4572 ;
  assign n13009 = n4547 | n4579 ;
  assign n13010 = x[93] & n4504 ;
  assign n13011 = n13009 | n13010 ;
  assign n13012 = n4672 | n13011 ;
  assign n30503 = ~n13012 ;
  assign n13013 = x[29] & n30503 ;
  assign n13014 = n28483 & n13012 ;
  assign n13015 = n13013 | n13014 ;
  assign n30504 = ~n13015 ;
  assign n13016 = n13008 & n30504 ;
  assign n30505 = ~n13008 ;
  assign n13671 = n30505 & n13015 ;
  assign n13672 = n13016 | n13671 ;
  assign n13673 = n13670 & n13672 ;
  assign n13694 = n13670 | n13672 ;
  assign n30506 = ~n13673 ;
  assign n13695 = n30506 & n13694 ;
  assign n30507 = ~n13693 ;
  assign n13696 = n30507 & n13695 ;
  assign n30508 = ~n13695 ;
  assign n14226 = n13693 & n30508 ;
  assign n14227 = n13696 | n14226 ;
  assign n14228 = n14225 & n14227 ;
  assign n14571 = n14225 | n14227 ;
  assign n30509 = ~n14228 ;
  assign n14572 = n30509 & n14571 ;
  assign n14573 = n14570 & n14572 ;
  assign n14575 = n14570 | n14572 ;
  assign n30510 = ~n14573 ;
  assign n14576 = n30510 & n14575 ;
  assign n15557 = n14620 | n15556 ;
  assign n15558 = n15516 & n15557 ;
  assign n15559 = n14586 | n15558 ;
  assign n30511 = ~n15559 ;
  assign n15560 = n14576 & n30511 ;
  assign n30512 = ~n14576 ;
  assign n15579 = n30512 & n15559 ;
  assign n15580 = n15560 | n15579 ;
  assign n7221 = n2867 & n7162 ;
  assign n7154 = x[100] & n7100 ;
  assign n7722 = x[101] & n7647 ;
  assign n15581 = n7154 | n7722 ;
  assign n15582 = x[102] & n7098 ;
  assign n15583 = n15581 | n15582 ;
  assign n15584 = n7221 | n15583 ;
  assign n30513 = ~n15584 ;
  assign n15585 = x[20] & n30513 ;
  assign n15586 = n28114 & n15584 ;
  assign n15587 = n15585 | n15586 ;
  assign n15588 = n15580 | n15587 ;
  assign n15589 = n15580 & n15587 ;
  assign n30514 = ~n15589 ;
  assign n16391 = n15588 & n30514 ;
  assign n30515 = ~n16218 ;
  assign n16392 = n30515 & n16391 ;
  assign n30516 = ~n16391 ;
  assign n16581 = n16218 & n30516 ;
  assign n16582 = n16392 | n16581 ;
  assign n16583 = n16578 | n16582 ;
  assign n16584 = n16578 & n16582 ;
  assign n30517 = ~n16584 ;
  assign n16585 = n16583 & n30517 ;
  assign n17440 = n16594 & n16597 ;
  assign n30518 = ~n16524 ;
  assign n16525 = n15608 & n30518 ;
  assign n30519 = ~n15608 ;
  assign n16586 = n30519 & n16524 ;
  assign n16587 = n16525 | n16586 ;
  assign n16595 = n16587 | n16594 ;
  assign n16596 = n16587 & n16594 ;
  assign n30520 = ~n16596 ;
  assign n17441 = n16595 & n30520 ;
  assign n17510 = n16611 | n17509 ;
  assign n17511 = n17441 & n17510 ;
  assign n17512 = n17440 | n17511 ;
  assign n30521 = ~n17512 ;
  assign n17513 = n16585 & n30521 ;
  assign n30522 = ~n16585 ;
  assign n17539 = n30522 & n17512 ;
  assign n17540 = n17513 | n17539 ;
  assign n10594 = n3876 & n10542 ;
  assign n10535 = x[106] & n10481 ;
  assign n11902 = x[107] & n11232 ;
  assign n17541 = n10535 | n11902 ;
  assign n17542 = x[108] & n10479 ;
  assign n17543 = n17541 | n17542 ;
  assign n17544 = n10594 | n17543 ;
  assign n30523 = ~n17544 ;
  assign n17545 = x[14] & n30523 ;
  assign n17546 = n27956 & n17544 ;
  assign n17547 = n17545 | n17546 ;
  assign n17548 = n17540 & n17547 ;
  assign n18258 = n17540 | n17547 ;
  assign n30524 = ~n17548 ;
  assign n18778 = n30524 & n18258 ;
  assign n30525 = ~n18778 ;
  assign n18779 = n18777 & n30525 ;
  assign n18259 = n18256 & n18258 ;
  assign n18260 = n17548 | n18259 ;
  assign n30526 = ~n18260 ;
  assign n18780 = n18258 & n30526 ;
  assign n18781 = n18779 | n18780 ;
  assign n12752 = n4246 & n12695 ;
  assign n12684 = x[109] & n12633 ;
  assign n14399 = x[110] & n13533 ;
  assign n18782 = n12684 | n14399 ;
  assign n18783 = x[111] & n12631 ;
  assign n18784 = n18782 | n18783 ;
  assign n18785 = n12752 | n18784 ;
  assign n30527 = ~n18785 ;
  assign n18786 = x[11] & n30527 ;
  assign n18787 = n27892 & n18785 ;
  assign n18788 = n18786 | n18787 ;
  assign n30528 = ~n18788 ;
  assign n18789 = n18781 & n30528 ;
  assign n30529 = ~n18781 ;
  assign n19557 = n30529 & n18788 ;
  assign n19558 = n18789 | n19557 ;
  assign n19559 = n19556 | n19558 ;
  assign n19560 = n19556 & n19558 ;
  assign n30530 = ~n19560 ;
  assign n20014 = n19559 & n30530 ;
  assign n30531 = ~n20013 ;
  assign n20015 = n30531 & n20014 ;
  assign n30532 = ~n20014 ;
  assign n20904 = n20013 & n30532 ;
  assign n20905 = n20015 | n20904 ;
  assign n20906 = n20903 | n20905 ;
  assign n20907 = n20903 & n20905 ;
  assign n30533 = ~n20907 ;
  assign n21047 = n20906 & n30533 ;
  assign n18418 = n797 & n18392 ;
  assign n18353 = x[115] & n18329 ;
  assign n18567 = x[116] & n18514 ;
  assign n21048 = n18353 | n18567 ;
  assign n21049 = x[117] & n18327 ;
  assign n21050 = n21048 | n21049 ;
  assign n21051 = n18418 | n21050 ;
  assign n30534 = ~n21051 ;
  assign n21052 = x[5] & n30534 ;
  assign n21053 = n27813 & n21051 ;
  assign n21054 = n21052 | n21053 ;
  assign n21055 = n21047 | n21054 ;
  assign n21056 = n21047 & n21054 ;
  assign n30535 = ~n21056 ;
  assign n22024 = n21055 & n30535 ;
  assign n22025 = n22023 & n22024 ;
  assign n22071 = n22023 | n22024 ;
  assign n30536 = ~n22025 ;
  assign n22072 = n30536 & n22071 ;
  assign n22073 = n22070 & n22072 ;
  assign n22074 = n22070 | n22072 ;
  assign n30537 = ~n22073 ;
  assign n22075 = n30537 & n22074 ;
  assign n23085 = n22085 | n23084 ;
  assign n23086 = n22075 & n23085 ;
  assign n27705 = n22075 | n23085 ;
  assign n30538 = ~n23086 ;
  assign n185 = n30538 & n27705 ;
  assign n22026 = n21056 | n22025 ;
  assign n18399 = n784 & n18392 ;
  assign n18386 = x[116] & n18329 ;
  assign n18564 = x[117] & n18514 ;
  assign n21035 = n18386 | n18564 ;
  assign n21036 = x[118] & n18327 ;
  assign n21037 = n21035 | n21036 ;
  assign n21038 = n18399 | n21037 ;
  assign n21039 = x[5] | n21038 ;
  assign n21040 = x[5] & n21038 ;
  assign n30539 = ~n21040 ;
  assign n21041 = n21039 & n30539 ;
  assign n20016 = n20013 & n20014 ;
  assign n20908 = n20016 | n20907 ;
  assign n15343 = n4474 & n15308 ;
  assign n15264 = x[113] & n15246 ;
  assign n17303 = x[114] & n16288 ;
  assign n19997 = n15264 | n17303 ;
  assign n19998 = x[115] & n15244 ;
  assign n19999 = n19997 | n19998 ;
  assign n20000 = n15343 | n19999 ;
  assign n30540 = ~n20000 ;
  assign n20001 = x[8] & n30540 ;
  assign n20002 = n27845 & n20000 ;
  assign n20003 = n20001 | n20002 ;
  assign n18790 = n18781 & n18788 ;
  assign n19561 = n18790 | n19560 ;
  assign n12747 = n4442 & n12695 ;
  assign n12662 = x[110] & n12633 ;
  assign n14375 = x[111] & n13533 ;
  assign n18674 = n12662 | n14375 ;
  assign n18675 = x[112] & n12631 ;
  assign n18676 = n18674 | n18675 ;
  assign n18677 = n12747 | n18676 ;
  assign n30541 = ~n18677 ;
  assign n18678 = x[11] & n30541 ;
  assign n18679 = n27892 & n18677 ;
  assign n18680 = n18678 | n18679 ;
  assign n10546 = n3639 & n10542 ;
  assign n10517 = x[107] & n10481 ;
  assign n11872 = x[108] & n11232 ;
  assign n17530 = n10517 | n11872 ;
  assign n17531 = x[109] & n10479 ;
  assign n17532 = n17530 | n17531 ;
  assign n17533 = n10546 | n17532 ;
  assign n30542 = ~n17533 ;
  assign n17534 = x[14] & n30542 ;
  assign n17535 = n27956 & n17533 ;
  assign n17536 = n17534 | n17535 ;
  assign n30543 = ~n14570 ;
  assign n14574 = n30543 & n14572 ;
  assign n30544 = ~n14572 ;
  assign n15514 = n14570 & n30544 ;
  assign n15515 = n14574 | n15514 ;
  assign n15561 = n15515 | n15559 ;
  assign n15562 = n15515 & n15559 ;
  assign n30545 = ~n15562 ;
  assign n15590 = n15561 & n30545 ;
  assign n30546 = ~n15587 ;
  assign n15591 = n30546 & n15590 ;
  assign n30547 = ~n15590 ;
  assign n15592 = n15587 & n30547 ;
  assign n15593 = n15591 | n15592 ;
  assign n16219 = n15593 | n16218 ;
  assign n16220 = n15593 & n16218 ;
  assign n30548 = ~n16220 ;
  assign n16571 = n16219 & n30548 ;
  assign n30549 = ~n16578 ;
  assign n16579 = n16571 & n30549 ;
  assign n30550 = ~n16571 ;
  assign n17438 = n30550 & n16578 ;
  assign n17439 = n16579 | n17438 ;
  assign n17514 = n17439 & n17512 ;
  assign n17515 = n16584 | n17514 ;
  assign n15563 = n14573 | n15562 ;
  assign n13697 = n13693 & n13695 ;
  assign n14229 = n13697 | n14228 ;
  assign n4664 = n2410 & n4632 ;
  assign n4531 = x[92] & n4514 ;
  assign n4604 = x[93] & n4572 ;
  assign n12995 = n4531 | n4604 ;
  assign n12996 = x[94] & n4504 ;
  assign n12997 = n12995 | n12996 ;
  assign n12998 = n4664 | n12997 ;
  assign n30551 = ~n12998 ;
  assign n12999 = x[29] & n30551 ;
  assign n13000 = n28483 & n12998 ;
  assign n13001 = n12999 | n13000 ;
  assign n12514 = n12512 & n12513 ;
  assign n12515 = n12107 | n12514 ;
  assign n10812 = n10803 & n10810 ;
  assign n11094 = n10812 | n11093 ;
  assign n3575 = n1239 & n3574 ;
  assign n3469 = x[83] & n3443 ;
  assign n3560 = x[84] & n3508 ;
  assign n10789 = n3469 | n3560 ;
  assign n10790 = x[85] & n3439 ;
  assign n10791 = n10789 | n10790 ;
  assign n10792 = n3575 | n10791 ;
  assign n30552 = ~n10792 ;
  assign n10793 = x[38] & n30552 ;
  assign n10794 = n28996 & n10792 ;
  assign n10795 = n10793 | n10794 ;
  assign n10093 = n10091 & n10092 ;
  assign n10329 = n10091 | n10092 ;
  assign n30553 = ~n10093 ;
  assign n10330 = n30553 & n10329 ;
  assign n10331 = n10327 & n10330 ;
  assign n10332 = n10093 | n10331 ;
  assign n3179 = n1003 & n3162 ;
  assign n3050 = x[80] & n3031 ;
  assign n3150 = x[81] & n3096 ;
  assign n10075 = n3050 | n3150 ;
  assign n10076 = x[82] & n3027 ;
  assign n10077 = n10075 | n10076 ;
  assign n10078 = n3179 | n10077 ;
  assign n30554 = ~n10078 ;
  assign n10079 = x[41] & n30554 ;
  assign n10080 = n29184 & n10078 ;
  assign n10081 = n10079 | n10080 ;
  assign n9447 = n9443 & n9445 ;
  assign n9637 = n9447 | n9636 ;
  assign n2641 = n1741 & n2635 ;
  assign n2508 = x[77] & n2492 ;
  assign n2564 = x[78] & n2557 ;
  assign n9427 = n2508 | n2564 ;
  assign n9428 = x[79] & n2488 ;
  assign n9429 = n9427 | n9428 ;
  assign n9430 = n2641 | n9429 ;
  assign n9431 = x[44] | n9430 ;
  assign n9432 = x[44] & n9430 ;
  assign n30555 = ~n9432 ;
  assign n9433 = n9431 & n30555 ;
  assign n8947 = n8943 & n8945 ;
  assign n9092 = n8947 | n9091 ;
  assign n2755 = n2321 & n2750 ;
  assign n2228 = x[74] & n2179 ;
  assign n2254 = x[75] & n2244 ;
  assign n8927 = n2228 | n2254 ;
  assign n8928 = x[76] & n2175 ;
  assign n8929 = n8927 | n8928 ;
  assign n8930 = n2755 | n8929 ;
  assign n30556 = ~n8930 ;
  assign n8931 = x[47] & n30556 ;
  assign n8932 = n29621 & n8930 ;
  assign n8933 = n8931 | n8932 ;
  assign n8451 = n8447 & n8449 ;
  assign n8452 = n8448 | n8451 ;
  assign n5985 = n1690 & n5976 ;
  assign n1577 = x[68] & n1551 ;
  assign n1642 = x[69] & n1616 ;
  assign n7883 = n1577 | n1642 ;
  assign n7884 = x[70] & n1547 ;
  assign n7885 = n7883 | n7884 ;
  assign n7886 = n5985 | n7885 ;
  assign n30557 = ~n7886 ;
  assign n7887 = x[53] & n30557 ;
  assign n7888 = n30125 & n7886 ;
  assign n7889 = n7887 | n7888 ;
  assign n27673 = x[56] & x[57] ;
  assign n1071 = x[56] | x[57] ;
  assign n30558 = ~n27673 ;
  assign n1072 = n30558 & n1071 ;
  assign n6849 = x[64] & n1072 ;
  assign n7417 = n7408 & n7415 ;
  assign n30559 = ~n6849 ;
  assign n7418 = n30559 & n7417 ;
  assign n30560 = ~n7417 ;
  assign n7420 = n6849 & n30560 ;
  assign n7421 = n7418 | n7420 ;
  assign n6506 = n1457 & n6494 ;
  assign n1370 = x[65] & n1319 ;
  assign n1403 = x[66] & n1384 ;
  assign n7422 = n1370 | n1403 ;
  assign n7423 = x[67] & n1315 ;
  assign n7424 = n7422 | n7423 ;
  assign n7425 = n6506 | n7424 ;
  assign n30561 = ~n7425 ;
  assign n7426 = x[56] & n30561 ;
  assign n7427 = n30379 & n7425 ;
  assign n7428 = n7426 | n7427 ;
  assign n7429 = n7421 | n7428 ;
  assign n7430 = n7421 & n7428 ;
  assign n30562 = ~n7430 ;
  assign n7890 = n7429 & n30562 ;
  assign n30563 = ~n7889 ;
  assign n7891 = n30563 & n7890 ;
  assign n30564 = ~n7890 ;
  assign n7957 = n7889 & n30564 ;
  assign n7958 = n7891 | n7957 ;
  assign n7959 = n7955 | n7958 ;
  assign n7960 = n7955 & n7958 ;
  assign n30565 = ~n7960 ;
  assign n8334 = n7959 & n30565 ;
  assign n3743 = n2007 & n3733 ;
  assign n1902 = x[71] & n1866 ;
  assign n1957 = x[72] & n1931 ;
  assign n8335 = n1902 | n1957 ;
  assign n8336 = x[73] & n1862 ;
  assign n8337 = n8335 | n8336 ;
  assign n8338 = n3743 | n8337 ;
  assign n30566 = ~n8338 ;
  assign n8339 = x[50] & n30566 ;
  assign n8340 = n29865 & n8338 ;
  assign n8341 = n8339 | n8340 ;
  assign n8342 = n8334 | n8341 ;
  assign n8343 = n8334 & n8341 ;
  assign n30567 = ~n8343 ;
  assign n8453 = n8342 & n30567 ;
  assign n8454 = n8452 & n8453 ;
  assign n8934 = n8452 | n8453 ;
  assign n30568 = ~n8454 ;
  assign n8935 = n30568 & n8934 ;
  assign n8936 = n8933 & n8935 ;
  assign n9093 = n8933 | n8935 ;
  assign n30569 = ~n8936 ;
  assign n9404 = n30569 & n9093 ;
  assign n30570 = ~n9092 ;
  assign n9406 = n30570 & n9404 ;
  assign n30571 = ~n9404 ;
  assign n9434 = n9092 & n30571 ;
  assign n9435 = n9406 | n9434 ;
  assign n9436 = n9433 & n9435 ;
  assign n9638 = n9433 | n9435 ;
  assign n30572 = ~n9436 ;
  assign n9639 = n30572 & n9638 ;
  assign n9640 = n9637 & n9639 ;
  assign n10082 = n9637 | n9639 ;
  assign n30573 = ~n9640 ;
  assign n10083 = n30573 & n10082 ;
  assign n30574 = ~n10081 ;
  assign n10333 = n30574 & n10083 ;
  assign n30575 = ~n10083 ;
  assign n10334 = n10081 & n30575 ;
  assign n10335 = n10333 | n10334 ;
  assign n10336 = n10332 & n10335 ;
  assign n10084 = n10081 & n10083 ;
  assign n30576 = ~n10084 ;
  assign n10796 = n10083 & n30576 ;
  assign n10797 = n10332 | n10796 ;
  assign n10798 = n10334 | n10797 ;
  assign n30577 = ~n10336 ;
  assign n10799 = n30577 & n10798 ;
  assign n10800 = n10795 | n10799 ;
  assign n10801 = n10795 & n10799 ;
  assign n30578 = ~n10801 ;
  assign n11095 = n10800 & n30578 ;
  assign n11096 = n11094 & n11095 ;
  assign n11354 = n11094 | n11095 ;
  assign n30579 = ~n11096 ;
  assign n11355 = n30579 & n11354 ;
  assign n4081 = n1720 & n4041 ;
  assign n3945 = x[86] & n3910 ;
  assign n4030 = x[87] & n3975 ;
  assign n11356 = n3945 | n4030 ;
  assign n11357 = x[88] & n3906 ;
  assign n11358 = n11356 | n11357 ;
  assign n11359 = n4081 | n11358 ;
  assign n30580 = ~n11359 ;
  assign n11360 = x[35] & n30580 ;
  assign n11361 = n28822 & n11359 ;
  assign n11362 = n11360 | n11361 ;
  assign n30581 = ~n11362 ;
  assign n11364 = n11355 & n30581 ;
  assign n30582 = ~n11355 ;
  assign n11365 = n30582 & n11362 ;
  assign n11366 = n11364 | n11365 ;
  assign n11697 = n11375 | n11696 ;
  assign n11698 = n11366 | n11697 ;
  assign n11699 = n11366 & n11697 ;
  assign n30583 = ~n11699 ;
  assign n12088 = n11698 & n30583 ;
  assign n2047 = n779 & n2046 ;
  assign n703 = x[89] & n663 ;
  assign n724 = x[90] & n720 ;
  assign n12089 = n703 | n724 ;
  assign n12090 = x[91] & n652 ;
  assign n12091 = n12089 | n12090 ;
  assign n12092 = n2047 | n12091 ;
  assign n30584 = ~n12092 ;
  assign n12093 = x[32] & n30584 ;
  assign n12094 = n28658 & n12092 ;
  assign n12095 = n12093 | n12094 ;
  assign n12096 = n12088 | n12095 ;
  assign n12097 = n12088 & n12095 ;
  assign n30585 = ~n12097 ;
  assign n12917 = n12096 & n30585 ;
  assign n30586 = ~n12515 ;
  assign n12919 = n30586 & n12917 ;
  assign n30587 = ~n12917 ;
  assign n13002 = n12515 & n30587 ;
  assign n13003 = n12919 | n13002 ;
  assign n13004 = n13001 & n13003 ;
  assign n13438 = n13001 | n13003 ;
  assign n30588 = ~n13004 ;
  assign n13439 = n30588 & n13438 ;
  assign n13017 = n13008 & n13015 ;
  assign n13674 = n13017 | n13673 ;
  assign n30589 = ~n13674 ;
  assign n13675 = n13439 & n30589 ;
  assign n30590 = ~n13439 ;
  assign n13676 = n30590 & n13674 ;
  assign n13677 = n13675 | n13676 ;
  assign n2440 = n452 & n2438 ;
  assign n373 = x[95] & n330 ;
  assign n392 = x[96] & n390 ;
  assign n13678 = n373 | n392 ;
  assign n13679 = x[97] & n322 ;
  assign n13680 = n13678 | n13679 ;
  assign n13681 = n2440 | n13680 ;
  assign n30591 = ~n13681 ;
  assign n13682 = x[26] & n30591 ;
  assign n13683 = n28342 & n13681 ;
  assign n13684 = n13682 | n13683 ;
  assign n30592 = ~n13684 ;
  assign n13685 = n13677 & n30592 ;
  assign n30593 = ~n13677 ;
  assign n14230 = n30593 & n13684 ;
  assign n14231 = n13685 | n14230 ;
  assign n14232 = n14229 | n14231 ;
  assign n14233 = n14229 & n14231 ;
  assign n30594 = ~n14233 ;
  assign n14554 = n14232 & n30594 ;
  assign n5310 = n2466 & n5302 ;
  assign n5270 = x[98] & n5240 ;
  assign n6279 = x[99] & n6179 ;
  assign n14555 = n5270 | n6279 ;
  assign n14556 = x[100] & n5238 ;
  assign n14557 = n14555 | n14556 ;
  assign n14558 = n5310 | n14557 ;
  assign n30595 = ~n14558 ;
  assign n14559 = x[23] & n30595 ;
  assign n14560 = n28221 & n14558 ;
  assign n14561 = n14559 | n14560 ;
  assign n14562 = n14554 | n14561 ;
  assign n14563 = n14554 & n14561 ;
  assign n30596 = ~n14563 ;
  assign n15564 = n14562 & n30596 ;
  assign n15565 = n15563 & n15564 ;
  assign n15566 = n15563 | n15564 ;
  assign n30597 = ~n15565 ;
  assign n15567 = n30597 & n15566 ;
  assign n7217 = n2626 & n7162 ;
  assign n7140 = x[101] & n7100 ;
  assign n7701 = x[102] & n7647 ;
  assign n15568 = n7140 | n7701 ;
  assign n15569 = x[103] & n7098 ;
  assign n15570 = n15568 | n15569 ;
  assign n15571 = n7217 | n15570 ;
  assign n30598 = ~n15571 ;
  assign n15572 = x[20] & n30598 ;
  assign n15573 = n28114 & n15571 ;
  assign n15574 = n15572 | n15573 ;
  assign n15576 = n15567 & n15574 ;
  assign n15577 = n15567 | n15574 ;
  assign n30599 = ~n15576 ;
  assign n15578 = n30599 & n15577 ;
  assign n16390 = n15587 & n15590 ;
  assign n16528 = n15607 | n16527 ;
  assign n16529 = n16391 & n16528 ;
  assign n16530 = n16390 | n16529 ;
  assign n30600 = ~n16530 ;
  assign n16531 = n15578 & n30600 ;
  assign n30601 = ~n15578 ;
  assign n16560 = n30601 & n16530 ;
  assign n16561 = n16531 | n16560 ;
  assign n8738 = n3223 & n8706 ;
  assign n8670 = x[104] & n8645 ;
  assign n9851 = x[105] & n9278 ;
  assign n16562 = n8670 | n9851 ;
  assign n16563 = x[106] & n8643 ;
  assign n16564 = n16562 | n16563 ;
  assign n16565 = n8738 | n16564 ;
  assign n30602 = ~n16565 ;
  assign n16566 = x[17] & n30602 ;
  assign n16567 = n28039 & n16565 ;
  assign n16568 = n16566 | n16567 ;
  assign n16569 = n16561 | n16568 ;
  assign n16570 = n16561 & n16568 ;
  assign n30603 = ~n16570 ;
  assign n17516 = n16569 & n30603 ;
  assign n17517 = n17515 & n17516 ;
  assign n17537 = n17515 | n17516 ;
  assign n30604 = ~n17517 ;
  assign n17538 = n30604 & n17537 ;
  assign n30605 = ~n17538 ;
  assign n18261 = n17536 & n30605 ;
  assign n30606 = ~n17536 ;
  assign n18262 = n30606 & n17538 ;
  assign n18263 = n18261 | n18262 ;
  assign n18264 = n18260 & n18263 ;
  assign n18681 = n18260 | n18262 ;
  assign n18682 = n18261 | n18681 ;
  assign n30607 = ~n18264 ;
  assign n18683 = n30607 & n18682 ;
  assign n30608 = ~n18683 ;
  assign n19562 = n18680 & n30608 ;
  assign n30609 = ~n18680 ;
  assign n19563 = n30609 & n18683 ;
  assign n19564 = n19562 | n19563 ;
  assign n19565 = n19561 & n19564 ;
  assign n20004 = n19561 | n19563 ;
  assign n20005 = n19562 | n20004 ;
  assign n30610 = ~n19565 ;
  assign n20006 = n30610 & n20005 ;
  assign n30611 = ~n20006 ;
  assign n20909 = n20003 & n30611 ;
  assign n30612 = ~n20003 ;
  assign n20910 = n30612 & n20006 ;
  assign n20911 = n20909 | n20910 ;
  assign n20912 = n20908 & n20911 ;
  assign n21042 = n20908 | n20910 ;
  assign n21043 = n20909 | n21042 ;
  assign n30613 = ~n20912 ;
  assign n21044 = n30613 & n21043 ;
  assign n30614 = ~n21044 ;
  assign n21045 = n21041 & n30614 ;
  assign n30615 = ~n21041 ;
  assign n22027 = n30615 & n21044 ;
  assign n22028 = n21045 | n22027 ;
  assign n22029 = n22026 | n22028 ;
  assign n22030 = n22026 & n22028 ;
  assign n30616 = ~n22030 ;
  assign n22052 = n22029 & n30616 ;
  assign n624 = n622 & n623 ;
  assign n625 = n23813 | n624 ;
  assign n27512 = x[120] & x[121] ;
  assign n626 = x[120] | x[121] ;
  assign n30617 = ~n27512 ;
  assign n4982 = n30617 & n626 ;
  assign n4983 = n625 | n4982 ;
  assign n4984 = n625 & n4982 ;
  assign n30618 = ~n4984 ;
  assign n4985 = n4983 & n30618 ;
  assign n19685 = n4985 & n19656 ;
  assign n19757 = x[119] & n19723 ;
  assign n19886 = x[120] & n19829 ;
  assign n22053 = n19757 | n19886 ;
  assign n22054 = x[121] & n19655 ;
  assign n22055 = n22053 | n22054 ;
  assign n22056 = n19685 | n22055 ;
  assign n30619 = ~n22056 ;
  assign n22057 = x[2] & n30619 ;
  assign n22058 = n27790 & n22056 ;
  assign n22059 = n22057 | n22058 ;
  assign n30620 = ~n22059 ;
  assign n22060 = n22052 & n30620 ;
  assign n30621 = ~n22052 ;
  assign n22062 = n30621 & n22059 ;
  assign n22063 = n22060 | n22062 ;
  assign n23087 = n22073 | n23086 ;
  assign n23088 = n22063 | n23087 ;
  assign n23089 = n22063 & n23087 ;
  assign n30622 = ~n23089 ;
  assign n186 = n23088 & n30622 ;
  assign n627 = n625 & n626 ;
  assign n628 = n27512 | n627 ;
  assign n23611 = x[121] & x[122] ;
  assign n629 = x[121] | x[122] ;
  assign n30623 = ~n23611 ;
  assign n5019 = n30623 & n629 ;
  assign n5020 = n628 & n5019 ;
  assign n5021 = n628 | n5019 ;
  assign n30624 = ~n5020 ;
  assign n5022 = n30624 & n5021 ;
  assign n19688 = n5022 & n19656 ;
  assign n19758 = x[120] & n19723 ;
  assign n19864 = x[121] & n19829 ;
  assign n22040 = n19758 | n19864 ;
  assign n22041 = x[122] & n19655 ;
  assign n22042 = n22040 | n22041 ;
  assign n22043 = n19688 | n22042 ;
  assign n22044 = x[2] | n22043 ;
  assign n22045 = x[2] & n22043 ;
  assign n30625 = ~n22045 ;
  assign n22046 = n22044 & n30625 ;
  assign n21046 = n21041 & n21044 ;
  assign n22031 = n21046 | n22030 ;
  assign n18419 = n5047 & n18392 ;
  assign n18379 = x[117] & n18329 ;
  assign n18548 = x[118] & n18514 ;
  assign n21025 = n18379 | n18548 ;
  assign n21026 = x[119] & n18327 ;
  assign n21027 = n21025 | n21026 ;
  assign n21028 = n18419 | n21027 ;
  assign n21029 = x[5] | n21028 ;
  assign n21030 = x[5] & n21028 ;
  assign n30626 = ~n21030 ;
  assign n21031 = n21029 & n30626 ;
  assign n20913 = n20003 & n20006 ;
  assign n20914 = n20912 | n20913 ;
  assign n15328 = n4702 & n15308 ;
  assign n15280 = x[114] & n15246 ;
  assign n17307 = x[115] & n16288 ;
  assign n19987 = n15280 | n17307 ;
  assign n19988 = x[116] & n15244 ;
  assign n19989 = n19987 | n19988 ;
  assign n19990 = n15328 | n19989 ;
  assign n19991 = x[8] | n19990 ;
  assign n19992 = x[8] & n19990 ;
  assign n30627 = ~n19992 ;
  assign n19993 = n19991 & n30627 ;
  assign n19566 = n18680 & n18683 ;
  assign n19567 = n19565 | n19566 ;
  assign n12755 = n4087 & n12695 ;
  assign n12681 = x[111] & n12633 ;
  assign n14352 = x[112] & n13533 ;
  assign n18664 = n12681 | n14352 ;
  assign n18665 = x[113] & n12631 ;
  assign n18666 = n18664 | n18665 ;
  assign n18667 = n12755 | n18666 ;
  assign n18668 = x[11] | n18667 ;
  assign n18669 = x[11] & n18667 ;
  assign n30628 = ~n18669 ;
  assign n18670 = n18668 & n30628 ;
  assign n18265 = n17536 & n17538 ;
  assign n18266 = n18264 | n18265 ;
  assign n13027 = n13018 & n13025 ;
  assign n13030 = n13025 | n13029 ;
  assign n30629 = ~n13031 ;
  assign n13032 = n13030 & n30629 ;
  assign n13431 = n13429 & n13430 ;
  assign n13432 = n13042 | n13431 ;
  assign n13433 = n13032 & n13432 ;
  assign n13434 = n13027 | n13433 ;
  assign n13435 = n13008 | n13015 ;
  assign n13436 = n13434 & n13435 ;
  assign n13437 = n13017 | n13436 ;
  assign n13440 = n13437 & n13439 ;
  assign n13441 = n13004 | n13440 ;
  assign n12918 = n12916 & n12917 ;
  assign n12920 = n12097 | n12918 ;
  assign n10337 = n10084 | n10336 ;
  assign n2728 = n2007 & n2722 ;
  assign n1896 = x[72] & n1866 ;
  assign n1959 = x[73] & n1931 ;
  assign n8321 = n1896 | n1959 ;
  assign n8322 = x[74] & n1862 ;
  assign n8323 = n8321 | n8322 ;
  assign n8324 = n2728 | n8323 ;
  assign n30630 = ~n8324 ;
  assign n8325 = x[50] & n30630 ;
  assign n8326 = n29865 & n8324 ;
  assign n8327 = n8325 | n8326 ;
  assign n7892 = n7889 & n7890 ;
  assign n7961 = n7892 | n7960 ;
  assign n4801 = n1690 & n4790 ;
  assign n1579 = x[69] & n1551 ;
  assign n1635 = x[70] & n1616 ;
  assign n7872 = n1579 | n1635 ;
  assign n7873 = x[71] & n1547 ;
  assign n7874 = n7872 | n7873 ;
  assign n7875 = n4801 | n7874 ;
  assign n30631 = ~n7875 ;
  assign n7876 = x[53] & n30631 ;
  assign n7877 = n30125 & n7875 ;
  assign n7878 = n7876 | n7877 ;
  assign n7419 = n6849 & n7417 ;
  assign n7431 = n7419 | n7430 ;
  assign n6418 = n1457 & n6408 ;
  assign n1347 = x[66] & n1319 ;
  assign n1408 = x[67] & n1384 ;
  assign n7387 = n1347 | n1408 ;
  assign n7388 = x[68] & n1315 ;
  assign n7389 = n7387 | n7388 ;
  assign n7390 = n6418 | n7389 ;
  assign n30632 = ~n7390 ;
  assign n7391 = x[56] & n30632 ;
  assign n7392 = n30379 & n7390 ;
  assign n7393 = n7391 | n7392 ;
  assign n6850 = x[59] & n30559 ;
  assign n27674 = x[58] & x[59] ;
  assign n1073 = x[58] | x[59] ;
  assign n30633 = ~n27674 ;
  assign n1074 = n30633 & n1073 ;
  assign n1217 = n1072 & n1074 ;
  assign n6449 = n1217 & n6437 ;
  assign n30634 = ~n1074 ;
  assign n1075 = n1072 & n30634 ;
  assign n6851 = x[65] & n1075 ;
  assign n27676 = x[57] & x[58] ;
  assign n1076 = x[57] | x[58] ;
  assign n30635 = ~n27676 ;
  assign n1077 = n30635 & n1076 ;
  assign n30636 = ~n1072 ;
  assign n1144 = n30636 & n1077 ;
  assign n6852 = x[64] & n1144 ;
  assign n6853 = n6851 | n6852 ;
  assign n6854 = n6449 | n6853 ;
  assign n30637 = ~n6854 ;
  assign n6855 = x[59] & n30637 ;
  assign n30638 = ~x[59] ;
  assign n6856 = n30638 & n6854 ;
  assign n6857 = n6855 | n6856 ;
  assign n30639 = ~n6857 ;
  assign n6858 = n6850 & n30639 ;
  assign n30640 = ~n6850 ;
  assign n7394 = n30640 & n6857 ;
  assign n7395 = n6858 | n7394 ;
  assign n30641 = ~n7393 ;
  assign n7396 = n30641 & n7395 ;
  assign n30642 = ~n7395 ;
  assign n7432 = n7393 & n30642 ;
  assign n7433 = n7396 | n7432 ;
  assign n30643 = ~n7431 ;
  assign n7434 = n30643 & n7433 ;
  assign n30644 = ~n7433 ;
  assign n7879 = n7431 & n30644 ;
  assign n7880 = n7434 | n7879 ;
  assign n30645 = ~n7878 ;
  assign n7881 = n30645 & n7880 ;
  assign n30646 = ~n7880 ;
  assign n7962 = n7878 & n30646 ;
  assign n7963 = n7881 | n7962 ;
  assign n7964 = n7961 & n7963 ;
  assign n8328 = n7961 | n7963 ;
  assign n30647 = ~n7964 ;
  assign n8329 = n30647 & n8328 ;
  assign n30648 = ~n8327 ;
  assign n8330 = n30648 & n8329 ;
  assign n30649 = ~n8329 ;
  assign n8332 = n8327 & n30649 ;
  assign n8333 = n8330 | n8332 ;
  assign n8455 = n8343 | n8454 ;
  assign n8456 = n8333 | n8455 ;
  assign n8457 = n8333 & n8455 ;
  assign n30650 = ~n8457 ;
  assign n8918 = n8456 & n30650 ;
  assign n2326 = n1775 & n2321 ;
  assign n2195 = x[75] & n2179 ;
  assign n2284 = x[76] & n2244 ;
  assign n8919 = n2195 | n2284 ;
  assign n8920 = x[77] & n2175 ;
  assign n8921 = n8919 | n8920 ;
  assign n8922 = n2326 | n8921 ;
  assign n30651 = ~n8922 ;
  assign n8923 = x[47] & n30651 ;
  assign n8924 = n29621 & n8922 ;
  assign n8925 = n8923 | n8924 ;
  assign n9096 = n8918 | n8925 ;
  assign n8926 = n8918 & n8925 ;
  assign n9094 = n9092 & n9093 ;
  assign n9095 = n8936 | n9094 ;
  assign n9097 = n9095 & n9096 ;
  assign n9099 = n8926 | n9097 ;
  assign n30652 = ~n9099 ;
  assign n9100 = n9096 & n30652 ;
  assign n30653 = ~n8926 ;
  assign n9098 = n30653 & n9096 ;
  assign n9405 = n9092 & n9404 ;
  assign n9407 = n8936 | n9405 ;
  assign n30654 = ~n9098 ;
  assign n9415 = n30654 & n9407 ;
  assign n9416 = n9100 | n9415 ;
  assign n2649 = n1270 & n2635 ;
  assign n2509 = x[78] & n2492 ;
  assign n2588 = x[79] & n2557 ;
  assign n9417 = n2509 | n2588 ;
  assign n9418 = x[80] & n2488 ;
  assign n9419 = n9417 | n9418 ;
  assign n9420 = n2649 | n9419 ;
  assign n30655 = ~n9420 ;
  assign n9421 = x[44] & n30655 ;
  assign n9422 = n29400 & n9420 ;
  assign n9423 = n9421 | n9422 ;
  assign n9424 = n9416 | n9423 ;
  assign n9425 = n9416 & n9423 ;
  assign n30656 = ~n9425 ;
  assign n9426 = n9424 & n30656 ;
  assign n9641 = n9436 | n9640 ;
  assign n30657 = ~n9641 ;
  assign n9642 = n9426 & n30657 ;
  assign n30658 = ~n9426 ;
  assign n10065 = n30658 & n9641 ;
  assign n10066 = n9642 | n10065 ;
  assign n3178 = n1057 & n3162 ;
  assign n3051 = x[81] & n3031 ;
  assign n3133 = x[82] & n3096 ;
  assign n10067 = n3051 | n3133 ;
  assign n10068 = x[83] & n3027 ;
  assign n10069 = n10067 | n10068 ;
  assign n10070 = n3178 | n10069 ;
  assign n30659 = ~n10070 ;
  assign n10071 = x[41] & n30659 ;
  assign n10072 = n29184 & n10070 ;
  assign n10073 = n10071 | n10072 ;
  assign n10074 = n10066 & n10073 ;
  assign n10338 = n10066 | n10073 ;
  assign n30660 = ~n10074 ;
  assign n10774 = n30660 & n10338 ;
  assign n30661 = ~n10774 ;
  assign n10775 = n10337 & n30661 ;
  assign n10751 = n10100 | n10102 ;
  assign n30662 = ~n10103 ;
  assign n10752 = n30662 & n10751 ;
  assign n10753 = n10308 & n10309 ;
  assign n10754 = n10140 | n10753 ;
  assign n10316 = n10125 & n10314 ;
  assign n10755 = n10125 | n10314 ;
  assign n30663 = ~n10316 ;
  assign n10756 = n30663 & n10755 ;
  assign n10757 = n10754 & n10756 ;
  assign n10758 = n10130 | n10757 ;
  assign n10759 = n10117 & n10758 ;
  assign n10760 = n10118 | n10759 ;
  assign n10761 = n10752 & n10760 ;
  assign n10762 = n10103 | n10761 ;
  assign n10766 = n10762 & n10764 ;
  assign n10767 = n10093 | n10766 ;
  assign n10768 = n10081 | n10083 ;
  assign n10769 = n30576 & n10768 ;
  assign n10770 = n10767 & n10769 ;
  assign n10771 = n10084 | n10770 ;
  assign n10772 = n10338 & n10771 ;
  assign n10773 = n10074 | n10772 ;
  assign n30664 = ~n10773 ;
  assign n10776 = n10338 & n30664 ;
  assign n10777 = n10775 | n10776 ;
  assign n3586 = n1213 & n3574 ;
  assign n3474 = x[84] & n3443 ;
  assign n3527 = x[85] & n3508 ;
  assign n10778 = n3474 | n3527 ;
  assign n10779 = x[86] & n3439 ;
  assign n10780 = n10778 | n10779 ;
  assign n10781 = n3586 | n10780 ;
  assign n30665 = ~n10781 ;
  assign n10782 = x[38] & n30665 ;
  assign n10783 = n28996 & n10781 ;
  assign n10784 = n10782 | n10783 ;
  assign n30666 = ~n10784 ;
  assign n10785 = n10777 & n30666 ;
  assign n30667 = ~n10777 ;
  assign n10787 = n30667 & n10784 ;
  assign n10788 = n10785 | n10787 ;
  assign n11097 = n10801 | n11096 ;
  assign n11098 = n10788 | n11097 ;
  assign n11099 = n10788 & n11097 ;
  assign n30668 = ~n11099 ;
  assign n11342 = n11098 & n30668 ;
  assign n4055 = n1453 & n4041 ;
  assign n3962 = x[87] & n3910 ;
  assign n4001 = x[88] & n3975 ;
  assign n11343 = n3962 | n4001 ;
  assign n11344 = x[89] & n3906 ;
  assign n11345 = n11343 | n11344 ;
  assign n11346 = n4055 | n11345 ;
  assign n30669 = ~n11346 ;
  assign n11347 = x[35] & n30669 ;
  assign n11348 = n28822 & n11346 ;
  assign n11349 = n11347 | n11348 ;
  assign n30670 = ~n11349 ;
  assign n11350 = n11342 & n30670 ;
  assign n30671 = ~n11342 ;
  assign n11352 = n30671 & n11349 ;
  assign n11353 = n11350 | n11352 ;
  assign n11363 = n11355 & n11362 ;
  assign n11700 = n11363 | n11699 ;
  assign n11701 = n11353 & n11700 ;
  assign n12077 = n11353 | n11700 ;
  assign n30672 = ~n11701 ;
  assign n12078 = n30672 & n12077 ;
  assign n1845 = n779 & n1841 ;
  assign n667 = x[90] & n663 ;
  assign n725 = x[91] & n720 ;
  assign n12079 = n667 | n725 ;
  assign n12080 = x[92] & n652 ;
  assign n12081 = n12079 | n12080 ;
  assign n12082 = n1845 | n12081 ;
  assign n30673 = ~n12082 ;
  assign n12083 = x[32] & n30673 ;
  assign n12084 = n28658 & n12082 ;
  assign n12085 = n12083 | n12084 ;
  assign n30674 = ~n12085 ;
  assign n12086 = n12078 & n30674 ;
  assign n30675 = ~n12078 ;
  assign n12921 = n30675 & n12085 ;
  assign n12922 = n12086 | n12921 ;
  assign n12923 = n12920 | n12922 ;
  assign n12924 = n12920 & n12922 ;
  assign n30676 = ~n12924 ;
  assign n12985 = n12923 & n30676 ;
  assign n4674 = n2152 & n4632 ;
  assign n4519 = x[93] & n4514 ;
  assign n4580 = x[94] & n4572 ;
  assign n12986 = n4519 | n4580 ;
  assign n12987 = x[95] & n4504 ;
  assign n12988 = n12986 | n12987 ;
  assign n12989 = n4674 | n12988 ;
  assign n30677 = ~n12989 ;
  assign n12990 = x[29] & n30677 ;
  assign n12991 = n28483 & n12989 ;
  assign n12992 = n12990 | n12991 ;
  assign n12993 = n12985 | n12992 ;
  assign n12994 = n12985 & n12992 ;
  assign n30678 = ~n12994 ;
  assign n13640 = n12993 & n30678 ;
  assign n13641 = n13441 | n13640 ;
  assign n13642 = n13441 & n13640 ;
  assign n30679 = ~n13642 ;
  assign n13643 = n13641 & n30679 ;
  assign n2843 = n452 & n2841 ;
  assign n387 = x[96] & n330 ;
  assign n396 = x[97] & n390 ;
  assign n13644 = n387 | n396 ;
  assign n13645 = x[98] & n322 ;
  assign n13646 = n13644 | n13645 ;
  assign n13647 = n2843 | n13646 ;
  assign n30680 = ~n13647 ;
  assign n13648 = x[26] & n30680 ;
  assign n13649 = n28342 & n13647 ;
  assign n13650 = n13648 | n13649 ;
  assign n30681 = ~n13650 ;
  assign n13651 = n13643 & n30681 ;
  assign n30682 = ~n13643 ;
  assign n13653 = n30682 & n13650 ;
  assign n13654 = n13651 | n13653 ;
  assign n13686 = n13677 & n13684 ;
  assign n14234 = n13686 | n14233 ;
  assign n14235 = n13654 & n14234 ;
  assign n14541 = n13654 | n14234 ;
  assign n30683 = ~n14235 ;
  assign n14542 = n30683 & n14541 ;
  assign n5336 = n2977 & n5302 ;
  assign n5287 = x[99] & n5240 ;
  assign n6261 = x[100] & n6179 ;
  assign n14543 = n5287 | n6261 ;
  assign n14544 = x[101] & n5238 ;
  assign n14545 = n14543 | n14544 ;
  assign n14546 = n5336 | n14545 ;
  assign n30684 = ~n14546 ;
  assign n14547 = x[23] & n30684 ;
  assign n14548 = n28221 & n14546 ;
  assign n14549 = n14547 | n14548 ;
  assign n30685 = ~n14549 ;
  assign n14550 = n14542 & n30685 ;
  assign n30686 = ~n14542 ;
  assign n14552 = n30686 & n14549 ;
  assign n14553 = n14550 | n14552 ;
  assign n15158 = n14586 | n15157 ;
  assign n15159 = n14576 & n15158 ;
  assign n15160 = n14573 | n15159 ;
  assign n15161 = n14562 & n15160 ;
  assign n15162 = n14563 | n15161 ;
  assign n15163 = n14553 & n15162 ;
  assign n15500 = n14553 | n15162 ;
  assign n30687 = ~n15163 ;
  assign n15501 = n30687 & n15500 ;
  assign n7216 = n3001 & n7162 ;
  assign n7156 = x[102] & n7100 ;
  assign n7717 = x[103] & n7647 ;
  assign n15502 = n7156 | n7717 ;
  assign n15503 = x[104] & n7098 ;
  assign n15504 = n15502 | n15503 ;
  assign n15505 = n7216 | n15504 ;
  assign n30688 = ~n15505 ;
  assign n15506 = x[20] & n30688 ;
  assign n15507 = n28114 & n15505 ;
  assign n15508 = n15506 | n15507 ;
  assign n30689 = ~n15508 ;
  assign n15511 = n15501 & n30689 ;
  assign n30690 = ~n15501 ;
  assign n15512 = n30690 & n15508 ;
  assign n15513 = n15511 | n15512 ;
  assign n16221 = n15589 | n16220 ;
  assign n16222 = n15578 & n16221 ;
  assign n16223 = n15576 | n16222 ;
  assign n16224 = n15513 | n16223 ;
  assign n16225 = n15513 & n16223 ;
  assign n30691 = ~n16225 ;
  assign n16551 = n16224 & n30691 ;
  assign n8762 = n3199 & n8706 ;
  assign n8694 = x[105] & n8645 ;
  assign n9855 = x[106] & n9278 ;
  assign n16552 = n8694 | n9855 ;
  assign n16553 = x[107] & n8643 ;
  assign n16554 = n16552 | n16553 ;
  assign n16555 = n8762 | n16554 ;
  assign n30692 = ~n16555 ;
  assign n16556 = x[17] & n30692 ;
  assign n16557 = n28039 & n16555 ;
  assign n16558 = n16556 | n16557 ;
  assign n17186 = n16551 | n16558 ;
  assign n16559 = n16551 & n16558 ;
  assign n16580 = n16571 & n16578 ;
  assign n17181 = n16596 | n17180 ;
  assign n17182 = n16585 & n17181 ;
  assign n17183 = n16580 | n17182 ;
  assign n17184 = n16569 & n17183 ;
  assign n17185 = n16570 | n17184 ;
  assign n17187 = n17185 & n17186 ;
  assign n17188 = n16559 | n17187 ;
  assign n30693 = ~n17188 ;
  assign n17189 = n17186 & n30693 ;
  assign n30694 = ~n16559 ;
  assign n17437 = n30694 & n17186 ;
  assign n17518 = n16570 | n17517 ;
  assign n30695 = ~n17437 ;
  assign n17519 = n30695 & n17518 ;
  assign n17520 = n17189 | n17519 ;
  assign n10598 = n3615 & n10542 ;
  assign n10532 = x[108] & n10481 ;
  assign n11903 = x[109] & n11232 ;
  assign n17521 = n10532 | n11903 ;
  assign n17522 = x[110] & n10479 ;
  assign n17523 = n17521 | n17522 ;
  assign n17524 = n10598 | n17523 ;
  assign n30696 = ~n17524 ;
  assign n17525 = x[14] & n30696 ;
  assign n17526 = n27956 & n17524 ;
  assign n17527 = n17525 | n17526 ;
  assign n17528 = n17520 | n17527 ;
  assign n17529 = n17520 & n17527 ;
  assign n30697 = ~n17529 ;
  assign n18267 = n17528 & n30697 ;
  assign n18268 = n18266 & n18267 ;
  assign n18671 = n18266 | n18267 ;
  assign n30698 = ~n18268 ;
  assign n18672 = n30698 & n18671 ;
  assign n18673 = n18670 & n18672 ;
  assign n19568 = n18670 | n18672 ;
  assign n30699 = ~n18673 ;
  assign n19569 = n30699 & n19568 ;
  assign n19570 = n19567 & n19569 ;
  assign n19994 = n19567 | n19569 ;
  assign n30700 = ~n19570 ;
  assign n19995 = n30700 & n19994 ;
  assign n19996 = n19993 & n19995 ;
  assign n20915 = n19993 | n19995 ;
  assign n30701 = ~n19996 ;
  assign n20916 = n30701 & n20915 ;
  assign n20917 = n20914 & n20916 ;
  assign n21032 = n20914 | n20916 ;
  assign n30702 = ~n20917 ;
  assign n21033 = n30702 & n21032 ;
  assign n21034 = n21031 & n21033 ;
  assign n22032 = n21031 | n21033 ;
  assign n30703 = ~n21034 ;
  assign n22033 = n30703 & n22032 ;
  assign n22034 = n22031 & n22033 ;
  assign n22047 = n22031 | n22033 ;
  assign n30704 = ~n22034 ;
  assign n22048 = n30704 & n22047 ;
  assign n22049 = n22046 & n22048 ;
  assign n22050 = n22046 | n22048 ;
  assign n30705 = ~n22049 ;
  assign n22051 = n30705 & n22050 ;
  assign n22061 = n22052 & n22059 ;
  assign n23090 = n22061 | n23089 ;
  assign n23091 = n22051 & n23090 ;
  assign n27708 = n22051 | n23090 ;
  assign n30706 = ~n23091 ;
  assign n187 = n30706 & n27708 ;
  assign n23092 = n22049 | n23091 ;
  assign n22035 = n21034 | n22034 ;
  assign n20918 = n19996 | n20917 ;
  assign n15339 = n797 & n15308 ;
  assign n15265 = x[115] & n15246 ;
  assign n17333 = x[116] & n16288 ;
  assign n19977 = n15265 | n17333 ;
  assign n19978 = x[117] & n15244 ;
  assign n19979 = n19977 | n19978 ;
  assign n19980 = n15339 | n19979 ;
  assign n30707 = ~n19980 ;
  assign n19981 = x[8] & n30707 ;
  assign n19982 = n27845 & n19980 ;
  assign n19983 = n19981 | n19982 ;
  assign n19571 = n18673 | n19570 ;
  assign n12738 = n4276 & n12695 ;
  assign n12680 = x[112] & n12633 ;
  assign n14385 = x[113] & n13533 ;
  assign n18654 = n12680 | n14385 ;
  assign n18655 = x[114] & n12631 ;
  assign n18656 = n18654 | n18655 ;
  assign n18657 = n12738 | n18656 ;
  assign n30708 = ~n18657 ;
  assign n18658 = x[11] & n30708 ;
  assign n18659 = n27892 & n18657 ;
  assign n18660 = n18658 | n18659 ;
  assign n18269 = n17529 | n18268 ;
  assign n15510 = n15501 & n15508 ;
  assign n16226 = n15510 | n16225 ;
  assign n2314 = n452 & n2313 ;
  assign n376 = x[97] & n330 ;
  assign n408 = x[98] & n390 ;
  assign n13627 = n376 | n408 ;
  assign n13628 = x[99] & n322 ;
  assign n13629 = n13627 | n13628 ;
  assign n13630 = n2314 | n13629 ;
  assign n30709 = ~n13630 ;
  assign n13631 = x[26] & n30709 ;
  assign n13632 = n28342 & n13630 ;
  assign n13633 = n13631 | n13632 ;
  assign n13442 = n12993 & n13441 ;
  assign n13443 = n12994 | n13442 ;
  assign n12087 = n12078 & n12085 ;
  assign n12925 = n12087 | n12924 ;
  assign n10786 = n10777 & n10784 ;
  assign n11100 = n10786 | n11099 ;
  assign n10339 = n10337 & n10338 ;
  assign n10340 = n10074 | n10339 ;
  assign n9643 = n9426 & n9641 ;
  assign n9644 = n9425 | n9643 ;
  assign n2661 = n1029 & n2635 ;
  assign n2541 = x[79] & n2492 ;
  assign n2616 = x[80] & n2557 ;
  assign n9397 = n2541 | n2616 ;
  assign n9398 = x[81] & n2488 ;
  assign n9399 = n9397 | n9398 ;
  assign n9400 = n2661 | n9399 ;
  assign n30710 = ~n9400 ;
  assign n9401 = x[44] & n30710 ;
  assign n9402 = n29400 & n9400 ;
  assign n9403 = n9401 | n9402 ;
  assign n2339 = n2084 & n2321 ;
  assign n2211 = x[76] & n2179 ;
  assign n2263 = x[77] & n2244 ;
  assign n8907 = n2211 | n2263 ;
  assign n8908 = x[78] & n2175 ;
  assign n8909 = n8907 | n8908 ;
  assign n8910 = n2339 | n8909 ;
  assign n30711 = ~n8910 ;
  assign n8911 = x[47] & n30711 ;
  assign n8912 = n29621 & n8910 ;
  assign n8913 = n8911 | n8912 ;
  assign n8331 = n8327 & n8329 ;
  assign n8458 = n8331 | n8457 ;
  assign n3295 = n2007 & n3289 ;
  assign n1899 = x[73] & n1866 ;
  assign n1961 = x[74] & n1931 ;
  assign n8310 = n1899 | n1961 ;
  assign n8311 = x[75] & n1862 ;
  assign n8312 = n8310 | n8311 ;
  assign n8313 = n3295 | n8312 ;
  assign n30712 = ~n8313 ;
  assign n8314 = x[50] & n30712 ;
  assign n8315 = n29865 & n8313 ;
  assign n8316 = n8314 | n8315 ;
  assign n7882 = n7878 & n7880 ;
  assign n7965 = n7882 | n7964 ;
  assign n7397 = n7393 & n7395 ;
  assign n7435 = n7431 & n7433 ;
  assign n7436 = n7397 | n7435 ;
  assign n6859 = n6850 & n6857 ;
  assign n6477 = n1217 & n6466 ;
  assign n1078 = n30636 & n1074 ;
  assign n30713 = ~n1077 ;
  assign n1079 = n30713 & n1078 ;
  assign n1116 = x[64] & n1079 ;
  assign n1193 = x[65] & n1144 ;
  assign n6860 = n1116 | n1193 ;
  assign n6861 = x[66] & n1075 ;
  assign n6862 = n6860 | n6861 ;
  assign n6863 = n6477 | n6862 ;
  assign n30714 = ~n6863 ;
  assign n6864 = x[59] & n30714 ;
  assign n6865 = n30638 & n6863 ;
  assign n6866 = n6864 | n6865 ;
  assign n30715 = ~n6866 ;
  assign n6867 = n6859 & n30715 ;
  assign n30716 = ~n6859 ;
  assign n7377 = n30716 & n6866 ;
  assign n7378 = n6867 | n7377 ;
  assign n6390 = n1457 & n6379 ;
  assign n1372 = x[67] & n1319 ;
  assign n1410 = x[68] & n1384 ;
  assign n7379 = n1372 | n1410 ;
  assign n7380 = x[69] & n1315 ;
  assign n7381 = n7379 | n7380 ;
  assign n7382 = n6390 | n7381 ;
  assign n30717 = ~n7382 ;
  assign n7383 = x[56] & n30717 ;
  assign n7384 = n30379 & n7382 ;
  assign n7385 = n7383 | n7384 ;
  assign n7386 = n7378 & n7385 ;
  assign n7437 = n7378 | n7385 ;
  assign n30718 = ~n7386 ;
  assign n7859 = n30718 & n7437 ;
  assign n30719 = ~n7859 ;
  assign n7860 = n7436 & n30719 ;
  assign n7438 = n7436 & n7437 ;
  assign n7439 = n7386 | n7438 ;
  assign n30720 = ~n7439 ;
  assign n7861 = n7437 & n30720 ;
  assign n7862 = n7860 | n7861 ;
  assign n3708 = n1690 & n3701 ;
  assign n1612 = x[70] & n1551 ;
  assign n1643 = x[71] & n1616 ;
  assign n7863 = n1612 | n1643 ;
  assign n7864 = x[72] & n1547 ;
  assign n7865 = n7863 | n7864 ;
  assign n7866 = n3708 | n7865 ;
  assign n30721 = ~n7866 ;
  assign n7867 = x[53] & n30721 ;
  assign n7868 = n30125 & n7866 ;
  assign n7869 = n7867 | n7868 ;
  assign n7870 = n7862 | n7869 ;
  assign n7871 = n7862 & n7869 ;
  assign n30722 = ~n7871 ;
  assign n7966 = n7870 & n30722 ;
  assign n30723 = ~n7965 ;
  assign n7967 = n30723 & n7966 ;
  assign n30724 = ~n7966 ;
  assign n8317 = n7965 & n30724 ;
  assign n8318 = n7967 | n8317 ;
  assign n30725 = ~n8316 ;
  assign n8319 = n30725 & n8318 ;
  assign n30726 = ~n8318 ;
  assign n8459 = n8316 & n30726 ;
  assign n8460 = n8319 | n8459 ;
  assign n30727 = ~n8458 ;
  assign n8461 = n30727 & n8460 ;
  assign n30728 = ~n8460 ;
  assign n8914 = n8458 & n30728 ;
  assign n8915 = n8461 | n8914 ;
  assign n8916 = n8913 | n8915 ;
  assign n8917 = n8913 & n8915 ;
  assign n30729 = ~n8917 ;
  assign n9101 = n8916 & n30729 ;
  assign n9408 = n9096 & n9407 ;
  assign n9409 = n8926 | n9408 ;
  assign n30730 = ~n9101 ;
  assign n9410 = n30730 & n9409 ;
  assign n30731 = ~n9409 ;
  assign n9411 = n9101 & n30731 ;
  assign n9412 = n9410 | n9411 ;
  assign n30732 = ~n9403 ;
  assign n9413 = n30732 & n9412 ;
  assign n30733 = ~n9412 ;
  assign n9645 = n9403 & n30733 ;
  assign n9646 = n9413 | n9645 ;
  assign n9647 = n9644 & n9646 ;
  assign n10054 = n9644 | n9646 ;
  assign n30734 = ~n9647 ;
  assign n10055 = n30734 & n10054 ;
  assign n3172 = n1293 & n3162 ;
  assign n3052 = x[82] & n3031 ;
  assign n3104 = x[83] & n3096 ;
  assign n10056 = n3052 | n3104 ;
  assign n10057 = x[84] & n3027 ;
  assign n10058 = n10056 | n10057 ;
  assign n10059 = n3172 | n10058 ;
  assign n30735 = ~n10059 ;
  assign n10060 = x[41] & n30735 ;
  assign n10061 = n29184 & n10059 ;
  assign n10062 = n10060 | n10061 ;
  assign n30736 = ~n10062 ;
  assign n10063 = n10055 & n30736 ;
  assign n30737 = ~n10055 ;
  assign n10341 = n30737 & n10062 ;
  assign n10342 = n10063 | n10341 ;
  assign n10343 = n10340 | n10342 ;
  assign n10344 = n10340 & n10342 ;
  assign n30738 = ~n10344 ;
  assign n10741 = n10343 & n30738 ;
  assign n3593 = n1522 & n3574 ;
  assign n3483 = x[85] & n3443 ;
  assign n3533 = x[86] & n3508 ;
  assign n10742 = n3483 | n3533 ;
  assign n10743 = x[87] & n3439 ;
  assign n10744 = n10742 | n10743 ;
  assign n10745 = n3593 | n10744 ;
  assign n30739 = ~n10745 ;
  assign n10746 = x[38] & n30739 ;
  assign n10747 = n28996 & n10745 ;
  assign n10748 = n10746 | n10747 ;
  assign n10749 = n10741 | n10748 ;
  assign n10750 = n10741 & n10748 ;
  assign n30740 = ~n10750 ;
  assign n11101 = n10749 & n30740 ;
  assign n11102 = n11100 & n11101 ;
  assign n11330 = n11100 | n11101 ;
  assign n30741 = ~n11102 ;
  assign n11331 = n30741 & n11330 ;
  assign n4077 = n1482 & n4041 ;
  assign n3964 = x[88] & n3910 ;
  assign n4032 = x[89] & n3975 ;
  assign n11332 = n3964 | n4032 ;
  assign n11333 = x[90] & n3906 ;
  assign n11334 = n11332 | n11333 ;
  assign n11335 = n4077 | n11334 ;
  assign n30742 = ~n11335 ;
  assign n11336 = x[35] & n30742 ;
  assign n11337 = n28822 & n11335 ;
  assign n11338 = n11336 | n11337 ;
  assign n11339 = n11331 | n11338 ;
  assign n11340 = n11331 & n11338 ;
  assign n30743 = ~n11340 ;
  assign n11341 = n11339 & n30743 ;
  assign n11351 = n11342 & n11349 ;
  assign n11702 = n11351 | n11701 ;
  assign n30744 = ~n11702 ;
  assign n11703 = n11341 & n30744 ;
  assign n30745 = ~n11341 ;
  assign n12067 = n30745 & n11702 ;
  assign n12068 = n11703 | n12067 ;
  assign n1688 = n779 & n1685 ;
  assign n670 = x[91] & n663 ;
  assign n726 = x[92] & n720 ;
  assign n12069 = n670 | n726 ;
  assign n12070 = x[93] & n652 ;
  assign n12071 = n12069 | n12070 ;
  assign n12072 = n1688 | n12071 ;
  assign n30746 = ~n12072 ;
  assign n12073 = x[32] & n30746 ;
  assign n12074 = n28658 & n12072 ;
  assign n12075 = n12073 | n12074 ;
  assign n12076 = n12068 & n12075 ;
  assign n12522 = n12068 | n12075 ;
  assign n30747 = ~n12076 ;
  assign n12972 = n30747 & n12522 ;
  assign n30748 = ~n12972 ;
  assign n12973 = n12925 & n30748 ;
  assign n12516 = n12096 & n12515 ;
  assign n12517 = n12097 | n12516 ;
  assign n12518 = n12078 | n12085 ;
  assign n30749 = ~n12087 ;
  assign n12519 = n30749 & n12518 ;
  assign n12520 = n12517 & n12519 ;
  assign n12521 = n12087 | n12520 ;
  assign n12523 = n12521 & n12522 ;
  assign n12524 = n12076 | n12523 ;
  assign n30750 = ~n12524 ;
  assign n12974 = n12522 & n30750 ;
  assign n12975 = n12973 | n12974 ;
  assign n4670 = n2000 & n4632 ;
  assign n4522 = x[94] & n4514 ;
  assign n4574 = x[95] & n4572 ;
  assign n12976 = n4522 | n4574 ;
  assign n12977 = x[96] & n4504 ;
  assign n12978 = n12976 | n12977 ;
  assign n12979 = n4670 | n12978 ;
  assign n30751 = ~n12979 ;
  assign n12980 = x[29] & n30751 ;
  assign n12981 = n28483 & n12979 ;
  assign n12982 = n12980 | n12981 ;
  assign n30752 = ~n12982 ;
  assign n12983 = n12975 & n30752 ;
  assign n30753 = ~n12975 ;
  assign n13444 = n30753 & n12982 ;
  assign n13445 = n12983 | n13444 ;
  assign n13446 = n13443 & n13445 ;
  assign n13634 = n13443 | n13445 ;
  assign n30754 = ~n13446 ;
  assign n13635 = n30754 & n13634 ;
  assign n30755 = ~n13633 ;
  assign n13636 = n30755 & n13635 ;
  assign n30756 = ~n13635 ;
  assign n13638 = n13633 & n30756 ;
  assign n13639 = n13636 | n13638 ;
  assign n13652 = n13643 & n13650 ;
  assign n14236 = n13652 | n14235 ;
  assign n30757 = ~n14236 ;
  assign n14237 = n13639 & n30757 ;
  assign n30758 = ~n13639 ;
  assign n14529 = n30758 & n14236 ;
  assign n14530 = n14237 | n14529 ;
  assign n5352 = n2867 & n5302 ;
  assign n5282 = x[100] & n5240 ;
  assign n6246 = x[101] & n6179 ;
  assign n14531 = n5282 | n6246 ;
  assign n14532 = x[102] & n5238 ;
  assign n14533 = n14531 | n14532 ;
  assign n14534 = n5352 | n14533 ;
  assign n30759 = ~n14534 ;
  assign n14535 = x[23] & n30759 ;
  assign n14536 = n28221 & n14534 ;
  assign n14537 = n14535 | n14536 ;
  assign n14538 = n14530 | n14537 ;
  assign n14539 = n14530 & n14537 ;
  assign n30760 = ~n14539 ;
  assign n14540 = n14538 & n30760 ;
  assign n14551 = n14542 & n14549 ;
  assign n15164 = n14551 | n15163 ;
  assign n30761 = ~n15164 ;
  assign n15165 = n14540 & n30761 ;
  assign n30762 = ~n14540 ;
  assign n15490 = n30762 & n15164 ;
  assign n15491 = n15165 | n15490 ;
  assign n7215 = n3409 & n7162 ;
  assign n7155 = x[103] & n7100 ;
  assign n7713 = x[104] & n7647 ;
  assign n15492 = n7155 | n7713 ;
  assign n15493 = x[105] & n7098 ;
  assign n15494 = n15492 | n15493 ;
  assign n15495 = n7215 | n15494 ;
  assign n30763 = ~n15495 ;
  assign n15496 = x[20] & n30763 ;
  assign n15497 = n28114 & n15495 ;
  assign n15498 = n15496 | n15497 ;
  assign n15499 = n15491 & n15498 ;
  assign n16227 = n15491 | n15498 ;
  assign n30764 = ~n15499 ;
  assign n16538 = n30764 & n16227 ;
  assign n30765 = ~n16538 ;
  assign n16539 = n16226 & n30765 ;
  assign n15509 = n15501 | n15508 ;
  assign n30766 = ~n15510 ;
  assign n16387 = n15509 & n30766 ;
  assign n30767 = ~n15574 ;
  assign n15575 = n15567 & n30767 ;
  assign n30768 = ~n15567 ;
  assign n16388 = n30768 & n15574 ;
  assign n16389 = n15575 | n16388 ;
  assign n16532 = n16389 & n16530 ;
  assign n16533 = n15576 | n16532 ;
  assign n16534 = n16387 & n16533 ;
  assign n16535 = n15510 | n16534 ;
  assign n16536 = n16227 & n16535 ;
  assign n16537 = n15499 | n16536 ;
  assign n30769 = ~n16537 ;
  assign n16540 = n16227 & n30769 ;
  assign n16541 = n16539 | n16540 ;
  assign n8765 = n3876 & n8706 ;
  assign n8687 = x[106] & n8645 ;
  assign n9869 = x[107] & n9278 ;
  assign n16542 = n8687 | n9869 ;
  assign n16543 = x[108] & n8643 ;
  assign n16544 = n16542 | n16543 ;
  assign n16545 = n8765 | n16544 ;
  assign n30770 = ~n16545 ;
  assign n16546 = x[17] & n30770 ;
  assign n16547 = n28039 & n16545 ;
  assign n16548 = n16546 | n16547 ;
  assign n30771 = ~n16548 ;
  assign n16549 = n16541 & n30771 ;
  assign n30772 = ~n16541 ;
  assign n17190 = n30772 & n16548 ;
  assign n17191 = n16549 | n17190 ;
  assign n17192 = n17188 | n17191 ;
  assign n17193 = n17188 & n17191 ;
  assign n30773 = ~n17193 ;
  assign n17427 = n17192 & n30773 ;
  assign n10558 = n4246 & n10542 ;
  assign n10531 = x[109] & n10481 ;
  assign n11890 = x[110] & n11232 ;
  assign n17428 = n10531 | n11890 ;
  assign n17429 = x[111] & n10479 ;
  assign n17430 = n17428 | n17429 ;
  assign n17431 = n10558 | n17430 ;
  assign n30774 = ~n17431 ;
  assign n17432 = x[14] & n30774 ;
  assign n17433 = n27956 & n17431 ;
  assign n17434 = n17432 | n17433 ;
  assign n17435 = n17427 | n17434 ;
  assign n17436 = n17427 & n17434 ;
  assign n30775 = ~n17436 ;
  assign n18270 = n17435 & n30775 ;
  assign n18271 = n18269 | n18270 ;
  assign n18272 = n18269 & n18270 ;
  assign n30776 = ~n18272 ;
  assign n18661 = n18271 & n30776 ;
  assign n30777 = ~n18660 ;
  assign n18662 = n30777 & n18661 ;
  assign n30778 = ~n18661 ;
  assign n19572 = n18660 & n30778 ;
  assign n19573 = n18662 | n19572 ;
  assign n19574 = n19571 | n19573 ;
  assign n19575 = n19571 & n19573 ;
  assign n30779 = ~n19575 ;
  assign n19984 = n19574 & n30779 ;
  assign n30780 = ~n19983 ;
  assign n19985 = n30780 & n19984 ;
  assign n30781 = ~n19984 ;
  assign n20919 = n19983 & n30781 ;
  assign n20920 = n19985 | n20919 ;
  assign n20921 = n20918 | n20920 ;
  assign n20922 = n20918 & n20920 ;
  assign n30782 = ~n20922 ;
  assign n21001 = n20921 & n30782 ;
  assign n18421 = n4678 & n18392 ;
  assign n18359 = x[118] & n18329 ;
  assign n18541 = x[119] & n18514 ;
  assign n21002 = n18359 | n18541 ;
  assign n21003 = x[120] & n18327 ;
  assign n21004 = n21002 | n21003 ;
  assign n21005 = n18421 | n21004 ;
  assign n30783 = ~n21005 ;
  assign n21006 = x[5] & n30783 ;
  assign n21007 = n27813 & n21005 ;
  assign n21008 = n21006 | n21007 ;
  assign n21009 = n21001 | n21008 ;
  assign n21010 = n21001 & n21008 ;
  assign n30784 = ~n21010 ;
  assign n21011 = n21009 & n30784 ;
  assign n630 = n628 & n629 ;
  assign n631 = n23611 | n630 ;
  assign n27470 = x[122] & x[123] ;
  assign n632 = x[122] | x[123] ;
  assign n30785 = ~n27470 ;
  assign n5414 = n30785 & n632 ;
  assign n5415 = n631 | n5414 ;
  assign n5416 = n631 & n5414 ;
  assign n30786 = ~n5416 ;
  assign n5417 = n5415 & n30786 ;
  assign n19698 = n5417 & n19656 ;
  assign n19755 = x[121] & n19723 ;
  assign n19871 = x[122] & n19829 ;
  assign n21012 = n19755 | n19871 ;
  assign n21013 = x[123] & n19655 ;
  assign n21014 = n21012 | n21013 ;
  assign n21015 = n19698 | n21014 ;
  assign n30787 = ~n21015 ;
  assign n21016 = x[2] & n30787 ;
  assign n21017 = n27790 & n21015 ;
  assign n21018 = n21016 | n21017 ;
  assign n30788 = ~n21018 ;
  assign n21019 = n21011 & n30788 ;
  assign n30789 = ~n21011 ;
  assign n22036 = n30789 & n21018 ;
  assign n22037 = n21019 | n22036 ;
  assign n22038 = n22035 | n22037 ;
  assign n22039 = n22035 & n22037 ;
  assign n30790 = ~n22039 ;
  assign n23093 = n22038 & n30790 ;
  assign n23094 = n23092 & n23093 ;
  assign n30791 = ~n22037 ;
  assign n27710 = n22035 & n30791 ;
  assign n30792 = ~n22035 ;
  assign n27711 = n30792 & n22037 ;
  assign n27712 = n23092 | n27711 ;
  assign n27713 = n27710 | n27712 ;
  assign n30793 = ~n23094 ;
  assign n188 = n30793 & n27713 ;
  assign n23095 = n22039 | n23094 ;
  assign n21020 = n21011 & n21018 ;
  assign n21021 = n21010 | n21020 ;
  assign n633 = n631 & n632 ;
  assign n634 = n27470 | n633 ;
  assign n23405 = x[123] & x[124] ;
  assign n635 = x[123] | x[124] ;
  assign n30794 = ~n23405 ;
  assign n5835 = n30794 & n635 ;
  assign n5836 = n634 & n5835 ;
  assign n5837 = n634 | n5835 ;
  assign n30795 = ~n5836 ;
  assign n5838 = n30795 & n5837 ;
  assign n19692 = n5838 & n19656 ;
  assign n19756 = x[122] & n19723 ;
  assign n19879 = x[123] & n19829 ;
  assign n20986 = n19756 | n19879 ;
  assign n20987 = x[124] & n19655 ;
  assign n20988 = n20986 | n20987 ;
  assign n20989 = n19692 | n20988 ;
  assign n20990 = x[2] | n20989 ;
  assign n20991 = x[2] & n20989 ;
  assign n30796 = ~n20991 ;
  assign n20992 = n20990 & n30796 ;
  assign n18422 = n4985 & n18392 ;
  assign n18357 = x[119] & n18329 ;
  assign n18538 = x[120] & n18514 ;
  assign n20976 = n18357 | n18538 ;
  assign n20977 = x[121] & n18327 ;
  assign n20978 = n20976 | n20977 ;
  assign n20979 = n18422 | n20978 ;
  assign n20980 = x[5] | n20979 ;
  assign n20981 = x[5] & n20979 ;
  assign n30797 = ~n20981 ;
  assign n20982 = n20980 & n30797 ;
  assign n19986 = n19983 & n19984 ;
  assign n20923 = n19986 | n20922 ;
  assign n15348 = n784 & n15308 ;
  assign n15273 = x[116] & n15246 ;
  assign n17317 = x[117] & n16288 ;
  assign n19965 = n15273 | n17317 ;
  assign n19966 = x[118] & n15244 ;
  assign n19967 = n19965 | n19966 ;
  assign n19968 = n15348 | n19967 ;
  assign n30798 = ~n19968 ;
  assign n19969 = x[8] & n30798 ;
  assign n19970 = n27845 & n19968 ;
  assign n19971 = n19969 | n19970 ;
  assign n18663 = n18660 & n18661 ;
  assign n19576 = n18663 | n19575 ;
  assign n12746 = n4474 & n12695 ;
  assign n12685 = x[113] & n12633 ;
  assign n14378 = x[114] & n13533 ;
  assign n18643 = n12685 | n14378 ;
  assign n18644 = x[115] & n12631 ;
  assign n18645 = n18643 | n18644 ;
  assign n18646 = n12746 | n18645 ;
  assign n30799 = ~n18646 ;
  assign n18647 = x[11] & n30799 ;
  assign n18648 = n27892 & n18646 ;
  assign n18649 = n18647 | n18648 ;
  assign n18273 = n17436 | n18272 ;
  assign n10596 = n4442 & n10542 ;
  assign n10528 = x[110] & n10481 ;
  assign n11894 = x[111] & n11232 ;
  assign n17416 = n10528 | n11894 ;
  assign n17417 = x[112] & n10479 ;
  assign n17418 = n17416 | n17417 ;
  assign n17419 = n10596 | n17418 ;
  assign n30800 = ~n17419 ;
  assign n17420 = x[14] & n30800 ;
  assign n17421 = n27956 & n17419 ;
  assign n17422 = n17420 | n17421 ;
  assign n16550 = n16541 & n16548 ;
  assign n17194 = n16550 | n17193 ;
  assign n8753 = n3639 & n8706 ;
  assign n8699 = x[107] & n8645 ;
  assign n9859 = x[108] & n9278 ;
  assign n16378 = n8699 | n9859 ;
  assign n16379 = x[109] & n8643 ;
  assign n16380 = n16378 | n16379 ;
  assign n16381 = n8753 | n16380 ;
  assign n30801 = ~n16381 ;
  assign n16382 = x[17] & n30801 ;
  assign n16383 = n28039 & n16381 ;
  assign n16384 = n16382 | n16383 ;
  assign n16228 = n16226 & n16227 ;
  assign n16229 = n15499 | n16228 ;
  assign n15166 = n14540 & n15164 ;
  assign n15167 = n14539 | n15166 ;
  assign n13637 = n13633 & n13635 ;
  assign n14238 = n13639 & n14236 ;
  assign n14239 = n13637 | n14238 ;
  assign n12984 = n12975 & n12982 ;
  assign n13447 = n12984 | n13446 ;
  assign n4669 = n2438 & n4632 ;
  assign n4541 = x[95] & n4514 ;
  assign n4586 = x[96] & n4572 ;
  assign n12961 = n4541 | n4586 ;
  assign n12962 = x[97] & n4504 ;
  assign n12963 = n12961 | n12962 ;
  assign n12964 = n4669 | n12963 ;
  assign n30802 = ~n12964 ;
  assign n12965 = x[29] & n30802 ;
  assign n12966 = n28483 & n12964 ;
  assign n12967 = n12965 | n12966 ;
  assign n10064 = n10055 & n10062 ;
  assign n10345 = n10064 | n10344 ;
  assign n3192 = n1239 & n3162 ;
  assign n3074 = x[83] & n3031 ;
  assign n3128 = x[84] & n3096 ;
  assign n10042 = n3074 | n3128 ;
  assign n10043 = x[85] & n3027 ;
  assign n10044 = n10042 | n10043 ;
  assign n10045 = n3192 | n10044 ;
  assign n30803 = ~n10045 ;
  assign n10046 = x[41] & n30803 ;
  assign n10047 = n29184 & n10045 ;
  assign n10048 = n10046 | n10047 ;
  assign n9414 = n9403 & n9412 ;
  assign n9648 = n9414 | n9647 ;
  assign n2644 = n1003 & n2635 ;
  assign n2554 = x[80] & n2492 ;
  assign n2565 = x[81] & n2557 ;
  assign n9387 = n2554 | n2565 ;
  assign n9388 = x[82] & n2488 ;
  assign n9389 = n9387 | n9388 ;
  assign n9390 = n2644 | n9389 ;
  assign n30804 = ~n9390 ;
  assign n9391 = x[44] & n30804 ;
  assign n9392 = n29400 & n9390 ;
  assign n9393 = n9391 | n9392 ;
  assign n9102 = n9099 & n9101 ;
  assign n9103 = n8917 | n9102 ;
  assign n2343 = n1741 & n2321 ;
  assign n2234 = x[77] & n2179 ;
  assign n2301 = x[78] & n2244 ;
  assign n8896 = n2234 | n2301 ;
  assign n8897 = x[79] & n2175 ;
  assign n8898 = n8896 | n8897 ;
  assign n8899 = n2343 | n8898 ;
  assign n30805 = ~n8899 ;
  assign n8900 = x[47] & n30805 ;
  assign n8901 = n29621 & n8899 ;
  assign n8902 = n8900 | n8901 ;
  assign n8320 = n8316 & n8318 ;
  assign n8462 = n8458 & n8460 ;
  assign n8463 = n8320 | n8462 ;
  assign n2753 = n2007 & n2750 ;
  assign n1903 = x[74] & n1866 ;
  assign n1934 = x[75] & n1931 ;
  assign n8299 = n1903 | n1934 ;
  assign n8300 = x[76] & n1862 ;
  assign n8301 = n8299 | n8300 ;
  assign n8302 = n2753 | n8301 ;
  assign n30806 = ~n8302 ;
  assign n8303 = x[50] & n30806 ;
  assign n8304 = n29865 & n8302 ;
  assign n8305 = n8303 | n8304 ;
  assign n7968 = n7965 & n7966 ;
  assign n7969 = n7871 | n7968 ;
  assign n5987 = n1457 & n5976 ;
  assign n1374 = x[68] & n1319 ;
  assign n1433 = x[69] & n1384 ;
  assign n7367 = n1374 | n1433 ;
  assign n7368 = x[70] & n1315 ;
  assign n7369 = n7367 | n7368 ;
  assign n7370 = n5987 | n7369 ;
  assign n30807 = ~n7370 ;
  assign n7371 = x[56] & n30807 ;
  assign n7372 = n30379 & n7370 ;
  assign n7373 = n7371 | n7372 ;
  assign n27665 = x[59] & x[60] ;
  assign n877 = x[59] | x[60] ;
  assign n30808 = ~n27665 ;
  assign n878 = n30808 & n877 ;
  assign n6431 = x[64] & n878 ;
  assign n6868 = n6859 & n6866 ;
  assign n30809 = ~n6431 ;
  assign n6869 = n30809 & n6868 ;
  assign n30810 = ~n6868 ;
  assign n6871 = n6431 & n30810 ;
  assign n6872 = n6869 | n6871 ;
  assign n6498 = n1217 & n6494 ;
  assign n1134 = x[65] & n1079 ;
  assign n1169 = x[66] & n1144 ;
  assign n6873 = n1134 | n1169 ;
  assign n6874 = x[67] & n1075 ;
  assign n6875 = n6873 | n6874 ;
  assign n6876 = n6498 | n6875 ;
  assign n30811 = ~n6876 ;
  assign n6877 = x[59] & n30811 ;
  assign n6878 = n30638 & n6876 ;
  assign n6879 = n6877 | n6878 ;
  assign n6880 = n6872 | n6879 ;
  assign n6881 = n6872 & n6879 ;
  assign n30812 = ~n6881 ;
  assign n7374 = n6880 & n30812 ;
  assign n30813 = ~n7373 ;
  assign n7375 = n30813 & n7374 ;
  assign n30814 = ~n7374 ;
  assign n7440 = n7373 & n30814 ;
  assign n7441 = n7375 | n7440 ;
  assign n7442 = n7439 | n7441 ;
  assign n7443 = n7439 & n7441 ;
  assign n30815 = ~n7443 ;
  assign n7849 = n7442 & n30815 ;
  assign n3739 = n1690 & n3733 ;
  assign n1599 = x[71] & n1551 ;
  assign n1664 = x[72] & n1616 ;
  assign n7850 = n1599 | n1664 ;
  assign n7851 = x[73] & n1547 ;
  assign n7852 = n7850 | n7851 ;
  assign n7853 = n3739 | n7852 ;
  assign n30816 = ~n7853 ;
  assign n7854 = x[53] & n30816 ;
  assign n7855 = n30125 & n7853 ;
  assign n7856 = n7854 | n7855 ;
  assign n7857 = n7849 | n7856 ;
  assign n7858 = n7849 & n7856 ;
  assign n30817 = ~n7858 ;
  assign n7970 = n7857 & n30817 ;
  assign n30818 = ~n7969 ;
  assign n7971 = n30818 & n7970 ;
  assign n30819 = ~n7970 ;
  assign n8306 = n7969 & n30819 ;
  assign n8307 = n7971 | n8306 ;
  assign n30820 = ~n8305 ;
  assign n8308 = n30820 & n8307 ;
  assign n30821 = ~n8307 ;
  assign n8464 = n8305 & n30821 ;
  assign n8465 = n8308 | n8464 ;
  assign n30822 = ~n8463 ;
  assign n8466 = n30822 & n8465 ;
  assign n30823 = ~n8465 ;
  assign n8903 = n8463 & n30823 ;
  assign n8904 = n8466 | n8903 ;
  assign n30824 = ~n8902 ;
  assign n8905 = n30824 & n8904 ;
  assign n30825 = ~n8904 ;
  assign n9104 = n8902 & n30825 ;
  assign n9105 = n8905 | n9104 ;
  assign n9106 = n9103 & n9105 ;
  assign n9394 = n9103 | n9105 ;
  assign n30826 = ~n9106 ;
  assign n9395 = n30826 & n9394 ;
  assign n30827 = ~n9395 ;
  assign n9649 = n9393 & n30827 ;
  assign n30828 = ~n9393 ;
  assign n9650 = n30828 & n9395 ;
  assign n9651 = n9649 | n9650 ;
  assign n9652 = n9648 & n9651 ;
  assign n10049 = n9648 | n9650 ;
  assign n10050 = n9649 | n10049 ;
  assign n30829 = ~n9652 ;
  assign n10051 = n30829 & n10050 ;
  assign n10052 = n10048 | n10051 ;
  assign n10053 = n10048 & n10051 ;
  assign n30830 = ~n10053 ;
  assign n10346 = n10052 & n30830 ;
  assign n10347 = n10345 & n10346 ;
  assign n10728 = n10345 | n10346 ;
  assign n30831 = ~n10347 ;
  assign n10729 = n30831 & n10728 ;
  assign n3591 = n1720 & n3574 ;
  assign n3489 = x[86] & n3443 ;
  assign n3531 = x[87] & n3508 ;
  assign n10730 = n3489 | n3531 ;
  assign n10731 = x[88] & n3439 ;
  assign n10732 = n10730 | n10731 ;
  assign n10733 = n3591 | n10732 ;
  assign n30832 = ~n10733 ;
  assign n10734 = x[38] & n30832 ;
  assign n10735 = n28996 & n10733 ;
  assign n10736 = n10734 | n10735 ;
  assign n30833 = ~n10736 ;
  assign n10737 = n10729 & n30833 ;
  assign n30834 = ~n10729 ;
  assign n10739 = n30834 & n10736 ;
  assign n10740 = n10737 | n10739 ;
  assign n11103 = n10750 | n11102 ;
  assign n11104 = n10740 | n11103 ;
  assign n11105 = n10740 & n11103 ;
  assign n30835 = ~n11105 ;
  assign n11318 = n11104 & n30835 ;
  assign n4060 = n2046 & n4041 ;
  assign n3969 = x[89] & n3910 ;
  assign n4036 = x[90] & n3975 ;
  assign n11319 = n3969 | n4036 ;
  assign n11320 = x[91] & n3906 ;
  assign n11321 = n11319 | n11320 ;
  assign n11322 = n4060 | n11321 ;
  assign n30836 = ~n11322 ;
  assign n11323 = x[35] & n30836 ;
  assign n11324 = n28822 & n11322 ;
  assign n11325 = n11323 | n11324 ;
  assign n30837 = ~n11325 ;
  assign n11327 = n11318 & n30837 ;
  assign n30838 = ~n11318 ;
  assign n11328 = n30838 & n11325 ;
  assign n11329 = n11327 | n11328 ;
  assign n11704 = n11341 & n11702 ;
  assign n11705 = n11340 | n11704 ;
  assign n11706 = n11329 | n11705 ;
  assign n11707 = n11329 & n11705 ;
  assign n30839 = ~n11707 ;
  assign n12058 = n11706 & n30839 ;
  assign n2411 = n779 & n2410 ;
  assign n674 = x[92] & n663 ;
  assign n748 = x[93] & n720 ;
  assign n12059 = n674 | n748 ;
  assign n12060 = x[94] & n652 ;
  assign n12061 = n12059 | n12060 ;
  assign n12062 = n2411 | n12061 ;
  assign n30840 = ~n12062 ;
  assign n12063 = x[32] & n30840 ;
  assign n12064 = n28658 & n12062 ;
  assign n12065 = n12063 | n12064 ;
  assign n12066 = n12058 & n12065 ;
  assign n12525 = n12058 | n12065 ;
  assign n30841 = ~n12066 ;
  assign n12526 = n30841 & n12525 ;
  assign n12926 = n12522 & n12925 ;
  assign n12927 = n12076 | n12926 ;
  assign n30842 = ~n12927 ;
  assign n12928 = n12526 & n30842 ;
  assign n30843 = ~n12526 ;
  assign n12968 = n30843 & n12927 ;
  assign n12969 = n12928 | n12968 ;
  assign n30844 = ~n12967 ;
  assign n12970 = n30844 & n12969 ;
  assign n30845 = ~n12969 ;
  assign n13448 = n12967 & n30845 ;
  assign n13449 = n12970 | n13448 ;
  assign n13450 = n13447 | n13449 ;
  assign n13451 = n13447 & n13449 ;
  assign n30846 = ~n13451 ;
  assign n13618 = n13450 & n30846 ;
  assign n2467 = n452 & n2466 ;
  assign n366 = x[98] & n330 ;
  assign n410 = x[99] & n390 ;
  assign n13619 = n366 | n410 ;
  assign n13620 = x[100] & n322 ;
  assign n13621 = n13619 | n13620 ;
  assign n13622 = n2467 | n13621 ;
  assign n30847 = ~n13622 ;
  assign n13623 = x[26] & n30847 ;
  assign n13624 = n28342 & n13622 ;
  assign n13625 = n13623 | n13624 ;
  assign n13626 = n13618 & n13625 ;
  assign n14240 = n13618 | n13625 ;
  assign n30848 = ~n13626 ;
  assign n14513 = n30848 & n14240 ;
  assign n30849 = ~n14239 ;
  assign n14514 = n30849 & n14513 ;
  assign n30850 = ~n14513 ;
  assign n14515 = n14239 & n30850 ;
  assign n14516 = n14514 | n14515 ;
  assign n5345 = n2626 & n5302 ;
  assign n5298 = x[101] & n5240 ;
  assign n6258 = x[102] & n6179 ;
  assign n14517 = n5298 | n6258 ;
  assign n14518 = x[103] & n5238 ;
  assign n14519 = n14517 | n14518 ;
  assign n14520 = n5345 | n14519 ;
  assign n30851 = ~n14520 ;
  assign n14521 = x[23] & n30851 ;
  assign n14522 = n28221 & n14520 ;
  assign n14523 = n14521 | n14522 ;
  assign n14524 = n14516 | n14523 ;
  assign n14525 = n14516 & n14523 ;
  assign n30852 = ~n14525 ;
  assign n15449 = n14524 & n30852 ;
  assign n30853 = ~n15167 ;
  assign n15450 = n30853 & n15449 ;
  assign n30854 = ~n15449 ;
  assign n15479 = n15167 & n30854 ;
  assign n15480 = n15450 | n15479 ;
  assign n7207 = n3223 & n7162 ;
  assign n7158 = x[104] & n7100 ;
  assign n7694 = x[105] & n7647 ;
  assign n15481 = n7158 | n7694 ;
  assign n15482 = x[106] & n7098 ;
  assign n15483 = n15481 | n15482 ;
  assign n15484 = n7207 | n15483 ;
  assign n30855 = ~n15484 ;
  assign n15485 = x[20] & n30855 ;
  assign n15486 = n28114 & n15484 ;
  assign n15487 = n15485 | n15486 ;
  assign n15488 = n15480 | n15487 ;
  assign n15489 = n15480 & n15487 ;
  assign n30856 = ~n15489 ;
  assign n16230 = n15488 & n30856 ;
  assign n30857 = ~n16229 ;
  assign n16231 = n30857 & n16230 ;
  assign n30858 = ~n16230 ;
  assign n16385 = n16229 & n30858 ;
  assign n16386 = n16231 | n16385 ;
  assign n30859 = ~n16386 ;
  assign n17195 = n16384 & n30859 ;
  assign n30860 = ~n16384 ;
  assign n17196 = n30860 & n16386 ;
  assign n17197 = n17195 | n17196 ;
  assign n17198 = n17194 & n17197 ;
  assign n17423 = n17194 | n17196 ;
  assign n17424 = n17195 | n17423 ;
  assign n30861 = ~n17198 ;
  assign n17425 = n30861 & n17424 ;
  assign n30862 = ~n17425 ;
  assign n18274 = n17422 & n30862 ;
  assign n30863 = ~n17422 ;
  assign n18275 = n30863 & n17425 ;
  assign n18276 = n18274 | n18275 ;
  assign n18277 = n18273 & n18276 ;
  assign n18650 = n18273 | n18275 ;
  assign n18651 = n18274 | n18650 ;
  assign n30864 = ~n18277 ;
  assign n18652 = n30864 & n18651 ;
  assign n30865 = ~n18652 ;
  assign n19577 = n18649 & n30865 ;
  assign n30866 = ~n18649 ;
  assign n19578 = n30866 & n18652 ;
  assign n19579 = n19577 | n19578 ;
  assign n19580 = n19576 & n19579 ;
  assign n19972 = n19576 | n19578 ;
  assign n19973 = n19577 | n19972 ;
  assign n30867 = ~n19580 ;
  assign n19974 = n30867 & n19973 ;
  assign n19975 = n19971 | n19974 ;
  assign n19976 = n19971 & n19974 ;
  assign n30868 = ~n19976 ;
  assign n20924 = n19975 & n30868 ;
  assign n20925 = n20923 & n20924 ;
  assign n20983 = n20923 | n20924 ;
  assign n30869 = ~n20925 ;
  assign n20984 = n30869 & n20983 ;
  assign n20985 = n20982 & n20984 ;
  assign n20993 = n20982 | n20984 ;
  assign n30870 = ~n20985 ;
  assign n20994 = n30870 & n20993 ;
  assign n20995 = n20992 & n20994 ;
  assign n21022 = n20992 | n20994 ;
  assign n30871 = ~n20995 ;
  assign n21023 = n30871 & n21022 ;
  assign n21024 = n21021 & n21023 ;
  assign n23096 = n21021 | n21023 ;
  assign n30872 = ~n21024 ;
  assign n23097 = n30872 & n23096 ;
  assign n23098 = n23095 & n23097 ;
  assign n27715 = n23095 | n23097 ;
  assign n30873 = ~n23098 ;
  assign n189 = n30873 & n27715 ;
  assign n15327 = n5047 & n15308 ;
  assign n15262 = x[117] & n15246 ;
  assign n17312 = x[118] & n16288 ;
  assign n19953 = n15262 | n17312 ;
  assign n19954 = x[119] & n15244 ;
  assign n19955 = n19953 | n19954 ;
  assign n19956 = n15327 | n19955 ;
  assign n19957 = x[8] | n19956 ;
  assign n19958 = x[8] & n19956 ;
  assign n30874 = ~n19958 ;
  assign n19959 = n19957 & n30874 ;
  assign n18653 = n18649 & n18652 ;
  assign n19581 = n18653 | n19580 ;
  assign n12740 = n4702 & n12695 ;
  assign n12660 = x[114] & n12633 ;
  assign n14374 = x[115] & n13533 ;
  assign n18633 = n12660 | n14374 ;
  assign n18634 = x[116] & n12631 ;
  assign n18635 = n18633 | n18634 ;
  assign n18636 = n12740 | n18635 ;
  assign n30875 = ~n18636 ;
  assign n18637 = x[11] & n30875 ;
  assign n18638 = n27892 & n18636 ;
  assign n18639 = n18637 | n18638 ;
  assign n17426 = n17422 & n17425 ;
  assign n18278 = n17426 | n18277 ;
  assign n10573 = n4087 & n10542 ;
  assign n10487 = x[111] & n10481 ;
  assign n11907 = x[112] & n11232 ;
  assign n17406 = n10487 | n11907 ;
  assign n17407 = x[113] & n10479 ;
  assign n17408 = n17406 | n17407 ;
  assign n17409 = n10573 | n17408 ;
  assign n17410 = x[14] | n17409 ;
  assign n17411 = x[14] & n17409 ;
  assign n30876 = ~n17411 ;
  assign n17412 = n17410 & n30876 ;
  assign n17199 = n16384 & n16386 ;
  assign n17200 = n17198 | n17199 ;
  assign n7199 = n3199 & n7162 ;
  assign n7147 = x[105] & n7100 ;
  assign n7674 = x[106] & n7647 ;
  assign n15471 = n7147 | n7674 ;
  assign n15472 = x[107] & n7098 ;
  assign n15473 = n15471 | n15472 ;
  assign n15474 = n7199 | n15473 ;
  assign n30877 = ~n15474 ;
  assign n15475 = x[20] & n30877 ;
  assign n15476 = n28114 & n15474 ;
  assign n15477 = n15475 | n15476 ;
  assign n12971 = n12967 & n12969 ;
  assign n13452 = n12971 | n13451 ;
  assign n12527 = n12524 & n12526 ;
  assign n12528 = n12066 | n12527 ;
  assign n8309 = n8305 & n8307 ;
  assign n8467 = n8463 & n8465 ;
  assign n8468 = n8309 | n8467 ;
  assign n2729 = n1690 & n2722 ;
  assign n1611 = x[72] & n1551 ;
  assign n1675 = x[73] & n1616 ;
  assign n7836 = n1611 | n1675 ;
  assign n7837 = x[74] & n1547 ;
  assign n7838 = n7836 | n7837 ;
  assign n7839 = n2729 | n7838 ;
  assign n30878 = ~n7839 ;
  assign n7840 = x[53] & n30878 ;
  assign n7841 = n30125 & n7839 ;
  assign n7842 = n7840 | n7841 ;
  assign n7376 = n7373 & n7374 ;
  assign n7444 = n7376 | n7443 ;
  assign n4799 = n1457 & n4790 ;
  assign n1358 = x[69] & n1319 ;
  assign n1424 = x[70] & n1384 ;
  assign n7356 = n1358 | n1424 ;
  assign n7357 = x[71] & n1315 ;
  assign n7358 = n7356 | n7357 ;
  assign n7359 = n4799 | n7358 ;
  assign n30879 = ~n7359 ;
  assign n7360 = x[56] & n30879 ;
  assign n7361 = n30379 & n7359 ;
  assign n7362 = n7360 | n7361 ;
  assign n6870 = n6431 & n6868 ;
  assign n6882 = n6870 | n6881 ;
  assign n6419 = n1217 & n6408 ;
  assign n1142 = x[66] & n1079 ;
  assign n1170 = x[67] & n1144 ;
  assign n6838 = n1142 | n1170 ;
  assign n6839 = x[68] & n1075 ;
  assign n6840 = n6838 | n6839 ;
  assign n6841 = n6419 | n6840 ;
  assign n30880 = ~n6841 ;
  assign n6842 = x[59] & n30880 ;
  assign n6843 = n30638 & n6841 ;
  assign n6844 = n6842 | n6843 ;
  assign n6432 = x[62] & n30809 ;
  assign n27667 = x[61] & x[62] ;
  assign n879 = x[61] | x[62] ;
  assign n30881 = ~n27667 ;
  assign n880 = n30881 & n879 ;
  assign n30882 = ~n880 ;
  assign n881 = n878 & n30882 ;
  assign n6433 = x[65] & n881 ;
  assign n27668 = x[60] & x[61] ;
  assign n897 = x[60] | x[61] ;
  assign n30883 = ~n27668 ;
  assign n898 = n30883 & n897 ;
  assign n30884 = ~n878 ;
  assign n949 = n30884 & n898 ;
  assign n6434 = x[64] & n949 ;
  assign n6435 = n6433 | n6434 ;
  assign n1006 = n878 & n880 ;
  assign n6450 = n1006 & n6437 ;
  assign n6452 = n6435 | n6450 ;
  assign n30885 = ~n6452 ;
  assign n6453 = x[62] & n30885 ;
  assign n30886 = ~x[62] ;
  assign n6454 = n30886 & n6452 ;
  assign n6455 = n6453 | n6454 ;
  assign n30887 = ~n6455 ;
  assign n6456 = n6432 & n30887 ;
  assign n30888 = ~n6432 ;
  assign n6845 = n30888 & n6455 ;
  assign n6846 = n6456 | n6845 ;
  assign n30889 = ~n6844 ;
  assign n6847 = n30889 & n6846 ;
  assign n30890 = ~n6846 ;
  assign n6883 = n6844 & n30890 ;
  assign n6884 = n6847 | n6883 ;
  assign n30891 = ~n6882 ;
  assign n6885 = n30891 & n6884 ;
  assign n30892 = ~n6884 ;
  assign n7363 = n6882 & n30892 ;
  assign n7364 = n6885 | n7363 ;
  assign n30893 = ~n7362 ;
  assign n7365 = n30893 & n7364 ;
  assign n30894 = ~n7364 ;
  assign n7445 = n7362 & n30894 ;
  assign n7446 = n7365 | n7445 ;
  assign n7447 = n7444 & n7446 ;
  assign n7843 = n7444 | n7446 ;
  assign n30895 = ~n7447 ;
  assign n7844 = n30895 & n7843 ;
  assign n30896 = ~n7842 ;
  assign n7845 = n30896 & n7844 ;
  assign n30897 = ~n7844 ;
  assign n7847 = n7842 & n30897 ;
  assign n7848 = n7845 | n7847 ;
  assign n7972 = n7969 & n7970 ;
  assign n7973 = n7858 | n7972 ;
  assign n7974 = n7848 | n7973 ;
  assign n7975 = n7848 & n7973 ;
  assign n30898 = ~n7975 ;
  assign n8290 = n7974 & n30898 ;
  assign n2017 = n1775 & n2007 ;
  assign n1914 = x[75] & n1866 ;
  assign n1990 = x[76] & n1931 ;
  assign n8291 = n1914 | n1990 ;
  assign n8292 = x[77] & n1862 ;
  assign n8293 = n8291 | n8292 ;
  assign n8294 = n2017 | n8293 ;
  assign n30899 = ~n8294 ;
  assign n8295 = x[50] & n30899 ;
  assign n8296 = n29865 & n8294 ;
  assign n8297 = n8295 | n8296 ;
  assign n8298 = n8290 & n8297 ;
  assign n8469 = n8290 | n8297 ;
  assign n30900 = ~n8298 ;
  assign n8470 = n30900 & n8469 ;
  assign n30901 = ~n8470 ;
  assign n8883 = n8468 & n30901 ;
  assign n8471 = n8468 & n8469 ;
  assign n8472 = n8298 | n8471 ;
  assign n30902 = ~n8472 ;
  assign n8884 = n8469 & n30902 ;
  assign n8885 = n8883 | n8884 ;
  assign n2335 = n1270 & n2321 ;
  assign n2205 = x[78] & n2179 ;
  assign n2305 = x[79] & n2244 ;
  assign n8886 = n2205 | n2305 ;
  assign n8887 = x[80] & n2175 ;
  assign n8888 = n8886 | n8887 ;
  assign n8889 = n2335 | n8888 ;
  assign n30903 = ~n8889 ;
  assign n8890 = x[47] & n30903 ;
  assign n8891 = n29621 & n8889 ;
  assign n8892 = n8890 | n8891 ;
  assign n8893 = n8885 | n8892 ;
  assign n8894 = n8885 & n8892 ;
  assign n30904 = ~n8894 ;
  assign n8895 = n8893 & n30904 ;
  assign n8906 = n8902 & n8904 ;
  assign n9107 = n8906 | n9106 ;
  assign n30905 = ~n9107 ;
  assign n9108 = n8895 & n30905 ;
  assign n30906 = ~n8895 ;
  assign n9377 = n30906 & n9107 ;
  assign n9378 = n9108 | n9377 ;
  assign n2642 = n1057 & n2635 ;
  assign n2531 = x[81] & n2492 ;
  assign n2614 = x[82] & n2557 ;
  assign n9379 = n2531 | n2614 ;
  assign n9380 = x[83] & n2488 ;
  assign n9381 = n9379 | n9380 ;
  assign n9382 = n2642 | n9381 ;
  assign n30907 = ~n9382 ;
  assign n9383 = x[44] & n30907 ;
  assign n9384 = n29400 & n9382 ;
  assign n9385 = n9383 | n9384 ;
  assign n9654 = n9378 | n9385 ;
  assign n9386 = n9378 & n9385 ;
  assign n9396 = n9393 & n9395 ;
  assign n9653 = n9396 | n9652 ;
  assign n9655 = n9653 & n9654 ;
  assign n9656 = n9386 | n9655 ;
  assign n30908 = ~n9656 ;
  assign n9657 = n9654 & n30908 ;
  assign n30909 = ~n9386 ;
  assign n10029 = n30909 & n9654 ;
  assign n30910 = ~n10029 ;
  assign n10030 = n9653 & n30910 ;
  assign n10031 = n9657 | n10030 ;
  assign n3191 = n1213 & n3162 ;
  assign n3091 = x[84] & n3031 ;
  assign n3146 = x[85] & n3096 ;
  assign n10032 = n3091 | n3146 ;
  assign n10033 = x[86] & n3027 ;
  assign n10034 = n10032 | n10033 ;
  assign n10035 = n3191 | n10034 ;
  assign n30911 = ~n10035 ;
  assign n10036 = x[41] & n30911 ;
  assign n10037 = n29184 & n10035 ;
  assign n10038 = n10036 | n10037 ;
  assign n10039 = n10031 | n10038 ;
  assign n10040 = n10031 & n10038 ;
  assign n30912 = ~n10040 ;
  assign n10041 = n10039 & n30912 ;
  assign n10348 = n10053 | n10347 ;
  assign n10349 = n10041 | n10348 ;
  assign n10350 = n10041 & n10348 ;
  assign n30913 = ~n10350 ;
  assign n10716 = n10349 & n30913 ;
  assign n3604 = n1453 & n3574 ;
  assign n3505 = x[87] & n3443 ;
  assign n3552 = x[88] & n3508 ;
  assign n10717 = n3505 | n3552 ;
  assign n10718 = x[89] & n3439 ;
  assign n10719 = n10717 | n10718 ;
  assign n10720 = n3604 | n10719 ;
  assign n30914 = ~n10720 ;
  assign n10721 = x[38] & n30914 ;
  assign n10722 = n28996 & n10720 ;
  assign n10723 = n10721 | n10722 ;
  assign n30915 = ~n10723 ;
  assign n10724 = n10716 & n30915 ;
  assign n30916 = ~n10716 ;
  assign n10726 = n30916 & n10723 ;
  assign n10727 = n10724 | n10726 ;
  assign n10738 = n10729 & n10736 ;
  assign n11106 = n10738 | n11105 ;
  assign n11107 = n10727 & n11106 ;
  assign n11305 = n10727 | n11106 ;
  assign n30917 = ~n11107 ;
  assign n11306 = n30917 & n11305 ;
  assign n4074 = n1841 & n4041 ;
  assign n3965 = x[90] & n3910 ;
  assign n4023 = x[91] & n3975 ;
  assign n11307 = n3965 | n4023 ;
  assign n11308 = x[92] & n3906 ;
  assign n11309 = n11307 | n11308 ;
  assign n11310 = n4074 | n11309 ;
  assign n30918 = ~n11310 ;
  assign n11311 = x[35] & n30918 ;
  assign n11312 = n28822 & n11310 ;
  assign n11313 = n11311 | n11312 ;
  assign n30919 = ~n11313 ;
  assign n11314 = n11306 & n30919 ;
  assign n30920 = ~n11306 ;
  assign n11316 = n30920 & n11313 ;
  assign n11317 = n11314 | n11316 ;
  assign n11326 = n11318 & n11325 ;
  assign n11708 = n11326 | n11707 ;
  assign n11709 = n11317 & n11708 ;
  assign n12047 = n11317 | n11708 ;
  assign n30921 = ~n11709 ;
  assign n12048 = n30921 & n12047 ;
  assign n2155 = n779 & n2152 ;
  assign n668 = x[93] & n663 ;
  assign n727 = x[94] & n720 ;
  assign n12049 = n668 | n727 ;
  assign n12050 = x[95] & n652 ;
  assign n12051 = n12049 | n12050 ;
  assign n12052 = n2155 | n12051 ;
  assign n30922 = ~n12052 ;
  assign n12053 = x[32] & n30922 ;
  assign n12054 = n28658 & n12052 ;
  assign n12055 = n12053 | n12054 ;
  assign n30923 = ~n12055 ;
  assign n12529 = n12048 & n30923 ;
  assign n30924 = ~n12048 ;
  assign n12530 = n30924 & n12055 ;
  assign n12531 = n12529 | n12530 ;
  assign n12532 = n12528 | n12531 ;
  assign n12533 = n12528 & n12531 ;
  assign n30925 = ~n12533 ;
  assign n12951 = n12532 & n30925 ;
  assign n4668 = n2841 & n4632 ;
  assign n4518 = x[96] & n4514 ;
  assign n4581 = x[97] & n4572 ;
  assign n12952 = n4518 | n4581 ;
  assign n12953 = x[98] & n4504 ;
  assign n12954 = n12952 | n12953 ;
  assign n12955 = n4668 | n12954 ;
  assign n30926 = ~n12955 ;
  assign n12956 = x[29] & n30926 ;
  assign n12957 = n28483 & n12955 ;
  assign n12958 = n12956 | n12957 ;
  assign n12959 = n12951 | n12958 ;
  assign n12960 = n12951 & n12958 ;
  assign n30927 = ~n12960 ;
  assign n13453 = n12959 & n30927 ;
  assign n13454 = n13452 & n13453 ;
  assign n13605 = n13452 | n13453 ;
  assign n30928 = ~n13454 ;
  assign n13606 = n30928 & n13605 ;
  assign n2979 = n452 & n2977 ;
  assign n379 = x[99] & n330 ;
  assign n419 = x[100] & n390 ;
  assign n13607 = n379 | n419 ;
  assign n13608 = x[101] & n322 ;
  assign n13609 = n13607 | n13608 ;
  assign n13610 = n2979 | n13609 ;
  assign n30929 = ~n13610 ;
  assign n13611 = x[26] & n30929 ;
  assign n13612 = n28342 & n13610 ;
  assign n13613 = n13611 | n13612 ;
  assign n30930 = ~n13613 ;
  assign n13614 = n13606 & n30930 ;
  assign n30931 = ~n13606 ;
  assign n13616 = n30931 & n13613 ;
  assign n13617 = n13614 | n13616 ;
  assign n14241 = n14239 & n14240 ;
  assign n14242 = n13626 | n14241 ;
  assign n14243 = n13617 & n14242 ;
  assign n14501 = n13617 | n14242 ;
  assign n30932 = ~n14243 ;
  assign n14502 = n30932 & n14501 ;
  assign n5335 = n3001 & n5302 ;
  assign n5296 = x[102] & n5240 ;
  assign n6244 = x[103] & n6179 ;
  assign n14503 = n5296 | n6244 ;
  assign n14504 = x[104] & n5238 ;
  assign n14505 = n14503 | n14504 ;
  assign n14506 = n5335 | n14505 ;
  assign n30933 = ~n14506 ;
  assign n14507 = x[23] & n30933 ;
  assign n14508 = n28221 & n14506 ;
  assign n14509 = n14507 | n14508 ;
  assign n14510 = n14502 | n14509 ;
  assign n14511 = n14502 & n14509 ;
  assign n30934 = ~n14511 ;
  assign n14512 = n14510 & n30934 ;
  assign n30935 = ~n14523 ;
  assign n14526 = n14516 & n30935 ;
  assign n30936 = ~n14516 ;
  assign n14527 = n30936 & n14523 ;
  assign n14528 = n14526 | n14527 ;
  assign n15168 = n14528 & n15167 ;
  assign n15169 = n14525 | n15168 ;
  assign n15170 = n14512 & n15169 ;
  assign n16359 = n14512 | n15169 ;
  assign n30937 = ~n15170 ;
  assign n16360 = n30937 & n16359 ;
  assign n16361 = n15477 | n16360 ;
  assign n16363 = n15477 & n16360 ;
  assign n16232 = n16229 & n16230 ;
  assign n16233 = n15489 | n16232 ;
  assign n16364 = n16233 & n16361 ;
  assign n16365 = n16363 | n16364 ;
  assign n30938 = ~n16365 ;
  assign n16366 = n16361 & n30938 ;
  assign n15451 = n15167 & n15449 ;
  assign n15452 = n14525 | n15451 ;
  assign n30939 = ~n15452 ;
  assign n15453 = n14512 & n30939 ;
  assign n30940 = ~n14512 ;
  assign n15469 = n30940 & n15452 ;
  assign n15470 = n15453 | n15469 ;
  assign n15478 = n15470 & n15477 ;
  assign n30941 = ~n15478 ;
  assign n16362 = n30941 & n16361 ;
  assign n30942 = ~n16362 ;
  assign n16367 = n16233 & n30942 ;
  assign n16368 = n16366 | n16367 ;
  assign n8764 = n3615 & n8706 ;
  assign n8678 = x[108] & n8645 ;
  assign n9862 = x[109] & n9278 ;
  assign n16369 = n8678 | n9862 ;
  assign n16370 = x[110] & n8643 ;
  assign n16371 = n16369 | n16370 ;
  assign n16372 = n8764 | n16371 ;
  assign n30943 = ~n16372 ;
  assign n16373 = x[17] & n30943 ;
  assign n16374 = n28039 & n16372 ;
  assign n16375 = n16373 | n16374 ;
  assign n16376 = n16368 | n16375 ;
  assign n16377 = n16368 & n16375 ;
  assign n30944 = ~n16377 ;
  assign n17201 = n16376 & n30944 ;
  assign n17202 = n17200 & n17201 ;
  assign n17413 = n17200 | n17201 ;
  assign n30945 = ~n17202 ;
  assign n17414 = n30945 & n17413 ;
  assign n17415 = n17412 & n17414 ;
  assign n18279 = n17412 | n17414 ;
  assign n30946 = ~n17415 ;
  assign n18280 = n30946 & n18279 ;
  assign n30947 = ~n18278 ;
  assign n18281 = n30947 & n18280 ;
  assign n30948 = ~n18280 ;
  assign n18640 = n18278 & n30948 ;
  assign n18641 = n18281 | n18640 ;
  assign n18642 = n18639 & n18641 ;
  assign n19582 = n18639 | n18641 ;
  assign n30949 = ~n18642 ;
  assign n19583 = n30949 & n19582 ;
  assign n19584 = n19581 & n19583 ;
  assign n19960 = n19581 | n19583 ;
  assign n30950 = ~n19584 ;
  assign n19961 = n30950 & n19960 ;
  assign n19962 = n19959 & n19961 ;
  assign n19963 = n19959 | n19961 ;
  assign n30951 = ~n19962 ;
  assign n19964 = n30951 & n19963 ;
  assign n20926 = n19976 | n20925 ;
  assign n30952 = ~n20926 ;
  assign n20927 = n19964 & n30952 ;
  assign n30953 = ~n19964 ;
  assign n20948 = n30953 & n20926 ;
  assign n20949 = n20927 | n20948 ;
  assign n18409 = n5022 & n18392 ;
  assign n18358 = x[120] & n18329 ;
  assign n18540 = x[121] & n18514 ;
  assign n20950 = n18358 | n18540 ;
  assign n20951 = x[122] & n18327 ;
  assign n20952 = n20950 | n20951 ;
  assign n20953 = n18409 | n20952 ;
  assign n30954 = ~n20953 ;
  assign n20954 = x[5] & n30954 ;
  assign n20955 = n27813 & n20953 ;
  assign n20956 = n20954 | n20955 ;
  assign n30955 = ~n20956 ;
  assign n20957 = n20949 & n30955 ;
  assign n30956 = ~n20949 ;
  assign n20959 = n30956 & n20956 ;
  assign n20960 = n20957 | n20959 ;
  assign n636 = n634 & n635 ;
  assign n637 = n23405 | n636 ;
  assign n27658 = x[124] & x[125] ;
  assign n638 = x[124] | x[125] ;
  assign n30957 = ~n27658 ;
  assign n639 = n30957 & n638 ;
  assign n30958 = ~n637 ;
  assign n640 = n30958 & n639 ;
  assign n30959 = ~n639 ;
  assign n641 = n637 & n30959 ;
  assign n642 = n640 | n641 ;
  assign n19697 = n642 & n19656 ;
  assign n19760 = x[123] & n19723 ;
  assign n19862 = x[124] & n19829 ;
  assign n20961 = n19760 | n19862 ;
  assign n20962 = x[125] & n19655 ;
  assign n20963 = n20961 | n20962 ;
  assign n20964 = n19697 | n20963 ;
  assign n30960 = ~n20964 ;
  assign n20965 = x[2] & n30960 ;
  assign n20966 = n27790 & n20964 ;
  assign n20967 = n20965 | n20966 ;
  assign n30961 = ~n20967 ;
  assign n20968 = n20960 & n30961 ;
  assign n30962 = ~n20960 ;
  assign n20974 = n30962 & n20967 ;
  assign n20975 = n20968 | n20974 ;
  assign n20996 = n20985 | n20995 ;
  assign n30963 = ~n20996 ;
  assign n20997 = n20975 & n30963 ;
  assign n30964 = ~n20975 ;
  assign n20999 = n30964 & n20996 ;
  assign n21000 = n20997 | n20999 ;
  assign n23099 = n21024 | n23098 ;
  assign n23100 = n21000 | n23099 ;
  assign n23101 = n21000 & n23099 ;
  assign n30965 = ~n23101 ;
  assign n190 = n23100 & n30965 ;
  assign n20998 = n20975 & n20996 ;
  assign n23102 = n20998 | n23101 ;
  assign n20958 = n20949 & n20956 ;
  assign n20969 = n20960 & n20967 ;
  assign n20970 = n20958 | n20969 ;
  assign n19585 = n18642 | n19584 ;
  assign n18282 = n18278 & n18280 ;
  assign n18283 = n17415 | n18282 ;
  assign n10595 = n4276 & n10542 ;
  assign n10513 = x[112] & n10481 ;
  assign n11897 = x[113] & n11232 ;
  assign n17394 = n10513 | n11897 ;
  assign n17395 = x[114] & n10479 ;
  assign n17396 = n17394 | n17395 ;
  assign n17397 = n10595 | n17396 ;
  assign n30966 = ~n17397 ;
  assign n17398 = x[14] & n30966 ;
  assign n17399 = n27956 & n17397 ;
  assign n17400 = n17398 | n17399 ;
  assign n17203 = n16377 | n17202 ;
  assign n16234 = n15470 | n15477 ;
  assign n16235 = n16233 & n16234 ;
  assign n16236 = n15478 | n16235 ;
  assign n15454 = n14512 & n15452 ;
  assign n15455 = n14511 | n15454 ;
  assign n12057 = n12048 & n12055 ;
  assign n12534 = n12057 | n12533 ;
  assign n10351 = n10040 | n10350 ;
  assign n9109 = n8895 & n9107 ;
  assign n9110 = n8894 | n9109 ;
  assign n2334 = n1029 & n2321 ;
  assign n2239 = x[79] & n2179 ;
  assign n2303 = x[80] & n2244 ;
  assign n8872 = n2239 | n2303 ;
  assign n8873 = x[81] & n2175 ;
  assign n8874 = n8872 | n8873 ;
  assign n8875 = n2334 | n8874 ;
  assign n30967 = ~n8875 ;
  assign n8876 = x[47] & n30967 ;
  assign n8877 = n29621 & n8875 ;
  assign n8878 = n8876 | n8877 ;
  assign n2085 = n2007 & n2084 ;
  assign n1918 = x[76] & n1866 ;
  assign n1987 = x[77] & n1931 ;
  assign n8279 = n1918 | n1987 ;
  assign n8280 = x[78] & n1862 ;
  assign n8281 = n8279 | n8280 ;
  assign n8282 = n2085 | n8281 ;
  assign n30968 = ~n8282 ;
  assign n8283 = x[50] & n30968 ;
  assign n8284 = n29865 & n8282 ;
  assign n8285 = n8283 | n8284 ;
  assign n7846 = n7842 & n7844 ;
  assign n7976 = n7846 | n7975 ;
  assign n3290 = n1690 & n3289 ;
  assign n1567 = x[73] & n1551 ;
  assign n1674 = x[74] & n1616 ;
  assign n7825 = n1567 | n1674 ;
  assign n7826 = x[75] & n1547 ;
  assign n7827 = n7825 | n7826 ;
  assign n7828 = n3290 | n7827 ;
  assign n30969 = ~n7828 ;
  assign n7829 = x[53] & n30969 ;
  assign n7830 = n30125 & n7828 ;
  assign n7831 = n7829 | n7830 ;
  assign n7366 = n7362 & n7364 ;
  assign n7448 = n7366 | n7447 ;
  assign n6848 = n6844 & n6846 ;
  assign n6886 = n6882 & n6884 ;
  assign n6887 = n6848 | n6886 ;
  assign n6457 = n6432 & n6455 ;
  assign n899 = n30884 & n880 ;
  assign n30970 = ~n898 ;
  assign n900 = n30970 & n899 ;
  assign n921 = x[64] & n900 ;
  assign n966 = x[65] & n949 ;
  assign n6458 = n921 | n966 ;
  assign n6459 = x[66] & n881 ;
  assign n6460 = n6458 | n6459 ;
  assign n6479 = n1006 & n6466 ;
  assign n6481 = n6460 | n6479 ;
  assign n30971 = ~n6481 ;
  assign n6482 = x[62] & n30971 ;
  assign n6483 = n30886 & n6481 ;
  assign n6484 = n6482 | n6483 ;
  assign n30972 = ~n6484 ;
  assign n6485 = n6457 & n30972 ;
  assign n30973 = ~n6457 ;
  assign n6828 = n30973 & n6484 ;
  assign n6829 = n6485 | n6828 ;
  assign n6391 = n1217 & n6379 ;
  assign n1101 = x[67] & n1079 ;
  assign n1178 = x[68] & n1144 ;
  assign n6830 = n1101 | n1178 ;
  assign n6831 = x[69] & n1075 ;
  assign n6832 = n6830 | n6831 ;
  assign n6833 = n6391 | n6832 ;
  assign n30974 = ~n6833 ;
  assign n6834 = x[59] & n30974 ;
  assign n6835 = n30638 & n6833 ;
  assign n6836 = n6834 | n6835 ;
  assign n6837 = n6829 & n6836 ;
  assign n6888 = n6829 | n6836 ;
  assign n30975 = ~n6837 ;
  assign n7344 = n30975 & n6888 ;
  assign n30976 = ~n7344 ;
  assign n7345 = n6887 & n30976 ;
  assign n6889 = n6887 & n6888 ;
  assign n6890 = n6837 | n6889 ;
  assign n30977 = ~n6890 ;
  assign n7346 = n6888 & n30977 ;
  assign n7347 = n7345 | n7346 ;
  assign n3705 = n1457 & n3701 ;
  assign n1348 = x[70] & n1319 ;
  assign n1422 = x[71] & n1384 ;
  assign n7348 = n1348 | n1422 ;
  assign n7349 = x[72] & n1315 ;
  assign n7350 = n7348 | n7349 ;
  assign n7351 = n3705 | n7350 ;
  assign n30978 = ~n7351 ;
  assign n7352 = x[56] & n30978 ;
  assign n7353 = n30379 & n7351 ;
  assign n7354 = n7352 | n7353 ;
  assign n7355 = n7347 | n7354 ;
  assign n7449 = n7347 & n7354 ;
  assign n30979 = ~n7449 ;
  assign n7450 = n7355 & n30979 ;
  assign n30980 = ~n7448 ;
  assign n7451 = n30980 & n7450 ;
  assign n30981 = ~n7450 ;
  assign n7832 = n7448 & n30981 ;
  assign n7833 = n7451 | n7832 ;
  assign n30982 = ~n7831 ;
  assign n7834 = n30982 & n7833 ;
  assign n30983 = ~n7833 ;
  assign n7977 = n7831 & n30983 ;
  assign n7978 = n7834 | n7977 ;
  assign n30984 = ~n7976 ;
  assign n7979 = n30984 & n7978 ;
  assign n30985 = ~n7978 ;
  assign n8286 = n7976 & n30985 ;
  assign n8287 = n7979 | n8286 ;
  assign n30986 = ~n8285 ;
  assign n8288 = n30986 & n8287 ;
  assign n30987 = ~n8287 ;
  assign n8473 = n8285 & n30987 ;
  assign n8474 = n8288 | n8473 ;
  assign n30988 = ~n8474 ;
  assign n8475 = n8472 & n30988 ;
  assign n8879 = n30902 & n8474 ;
  assign n8880 = n8475 | n8879 ;
  assign n30989 = ~n8878 ;
  assign n8881 = n30989 & n8880 ;
  assign n30990 = ~n8880 ;
  assign n9111 = n8878 & n30990 ;
  assign n9112 = n8881 | n9111 ;
  assign n30991 = ~n9112 ;
  assign n9113 = n9110 & n30991 ;
  assign n30992 = ~n9110 ;
  assign n9366 = n30992 & n9112 ;
  assign n9367 = n9113 | n9366 ;
  assign n2658 = n1293 & n2635 ;
  assign n2553 = x[82] & n2492 ;
  assign n2601 = x[83] & n2557 ;
  assign n9368 = n2553 | n2601 ;
  assign n9369 = x[84] & n2488 ;
  assign n9370 = n9368 | n9369 ;
  assign n9371 = n2658 | n9370 ;
  assign n30993 = ~n9371 ;
  assign n9372 = x[44] & n30993 ;
  assign n9373 = n29400 & n9371 ;
  assign n9374 = n9372 | n9373 ;
  assign n30994 = ~n9374 ;
  assign n9375 = n9367 & n30994 ;
  assign n30995 = ~n9367 ;
  assign n9658 = n30995 & n9374 ;
  assign n9659 = n9375 | n9658 ;
  assign n9660 = n9656 | n9659 ;
  assign n9661 = n9656 & n9659 ;
  assign n30996 = ~n9661 ;
  assign n10019 = n9660 & n30996 ;
  assign n3187 = n1522 & n3162 ;
  assign n3068 = x[85] & n3031 ;
  assign n3154 = x[86] & n3096 ;
  assign n10020 = n3068 | n3154 ;
  assign n10021 = x[87] & n3027 ;
  assign n10022 = n10020 | n10021 ;
  assign n10023 = n3187 | n10022 ;
  assign n30997 = ~n10023 ;
  assign n10024 = x[41] & n30997 ;
  assign n10025 = n29184 & n10023 ;
  assign n10026 = n10024 | n10025 ;
  assign n10027 = n10019 | n10026 ;
  assign n10028 = n10019 & n10026 ;
  assign n30998 = ~n10028 ;
  assign n10352 = n10027 & n30998 ;
  assign n10353 = n10351 & n10352 ;
  assign n10703 = n10351 | n10352 ;
  assign n30999 = ~n10353 ;
  assign n10704 = n30999 & n10703 ;
  assign n3597 = n1482 & n3574 ;
  assign n3453 = x[88] & n3443 ;
  assign n3519 = x[89] & n3508 ;
  assign n10705 = n3453 | n3519 ;
  assign n10706 = x[90] & n3439 ;
  assign n10707 = n10705 | n10706 ;
  assign n10708 = n3597 | n10707 ;
  assign n31000 = ~n10708 ;
  assign n10709 = x[38] & n31000 ;
  assign n10710 = n28996 & n10708 ;
  assign n10711 = n10709 | n10710 ;
  assign n31001 = ~n10711 ;
  assign n10712 = n10704 & n31001 ;
  assign n31002 = ~n10704 ;
  assign n10714 = n31002 & n10711 ;
  assign n10715 = n10712 | n10714 ;
  assign n10725 = n10716 & n10723 ;
  assign n11108 = n10725 | n11107 ;
  assign n31003 = ~n11108 ;
  assign n11109 = n10715 & n31003 ;
  assign n31004 = ~n10715 ;
  assign n11292 = n31004 & n11108 ;
  assign n11293 = n11109 | n11292 ;
  assign n4080 = n1685 & n4041 ;
  assign n3938 = x[91] & n3910 ;
  assign n4022 = x[92] & n3975 ;
  assign n11294 = n3938 | n4022 ;
  assign n11295 = x[93] & n3906 ;
  assign n11296 = n11294 | n11295 ;
  assign n11297 = n4080 | n11296 ;
  assign n31005 = ~n11297 ;
  assign n11298 = x[35] & n31005 ;
  assign n11299 = n28822 & n11297 ;
  assign n11300 = n11298 | n11299 ;
  assign n31006 = ~n11300 ;
  assign n11301 = n11293 & n31006 ;
  assign n31007 = ~n11293 ;
  assign n11303 = n31007 & n11300 ;
  assign n11304 = n11301 | n11303 ;
  assign n11315 = n11306 & n11313 ;
  assign n11710 = n11315 | n11709 ;
  assign n31008 = ~n11710 ;
  assign n11711 = n11304 & n31008 ;
  assign n31009 = ~n11304 ;
  assign n12037 = n31009 & n11710 ;
  assign n12038 = n11711 | n12037 ;
  assign n2002 = n779 & n2000 ;
  assign n680 = x[94] & n663 ;
  assign n738 = x[95] & n720 ;
  assign n12039 = n680 | n738 ;
  assign n12040 = x[96] & n652 ;
  assign n12041 = n12039 | n12040 ;
  assign n12042 = n2002 | n12041 ;
  assign n31010 = ~n12042 ;
  assign n12043 = x[32] & n31010 ;
  assign n12044 = n28658 & n12042 ;
  assign n12045 = n12043 | n12044 ;
  assign n12046 = n12038 & n12045 ;
  assign n12535 = n12038 | n12045 ;
  assign n31011 = ~n12046 ;
  assign n12936 = n31011 & n12535 ;
  assign n31012 = ~n12936 ;
  assign n12937 = n12534 & n31012 ;
  assign n12929 = n12525 & n12927 ;
  assign n12930 = n12066 | n12929 ;
  assign n12056 = n12048 | n12055 ;
  assign n31013 = ~n12057 ;
  assign n12931 = n12056 & n31013 ;
  assign n12932 = n12930 & n12931 ;
  assign n12933 = n12057 | n12932 ;
  assign n12934 = n12535 & n12933 ;
  assign n12935 = n12046 | n12934 ;
  assign n31014 = ~n12935 ;
  assign n12938 = n12535 & n31014 ;
  assign n12939 = n12937 | n12938 ;
  assign n4666 = n2313 & n4632 ;
  assign n4517 = x[97] & n4514 ;
  assign n4583 = x[98] & n4572 ;
  assign n12940 = n4517 | n4583 ;
  assign n12941 = x[99] & n4504 ;
  assign n12942 = n12940 | n12941 ;
  assign n12943 = n4666 | n12942 ;
  assign n31015 = ~n12943 ;
  assign n12944 = x[29] & n31015 ;
  assign n12945 = n28483 & n12943 ;
  assign n12946 = n12944 | n12945 ;
  assign n31016 = ~n12946 ;
  assign n12947 = n12939 & n31016 ;
  assign n31017 = ~n12939 ;
  assign n12949 = n31017 & n12946 ;
  assign n12950 = n12947 | n12949 ;
  assign n13455 = n12960 | n13454 ;
  assign n13456 = n12950 & n13455 ;
  assign n13593 = n12950 | n13455 ;
  assign n31018 = ~n13456 ;
  assign n13594 = n31018 & n13593 ;
  assign n2868 = n452 & n2867 ;
  assign n351 = x[100] & n330 ;
  assign n393 = x[101] & n390 ;
  assign n13595 = n351 | n393 ;
  assign n13596 = x[102] & n322 ;
  assign n13597 = n13595 | n13596 ;
  assign n13598 = n2868 | n13597 ;
  assign n31019 = ~n13598 ;
  assign n13599 = x[26] & n31019 ;
  assign n13600 = n28342 & n13598 ;
  assign n13601 = n13599 | n13600 ;
  assign n13602 = n13594 | n13601 ;
  assign n13603 = n13594 & n13601 ;
  assign n31020 = ~n13603 ;
  assign n13604 = n13602 & n31020 ;
  assign n13615 = n13606 & n13613 ;
  assign n14244 = n13615 | n14243 ;
  assign n14245 = n13604 | n14244 ;
  assign n14246 = n13604 & n14244 ;
  assign n31021 = ~n14246 ;
  assign n14492 = n14245 & n31021 ;
  assign n5338 = n3409 & n5302 ;
  assign n5266 = x[103] & n5240 ;
  assign n6264 = x[104] & n6179 ;
  assign n14493 = n5266 | n6264 ;
  assign n14494 = x[105] & n5238 ;
  assign n14495 = n14493 | n14494 ;
  assign n14496 = n5338 | n14495 ;
  assign n31022 = ~n14496 ;
  assign n14497 = x[23] & n31022 ;
  assign n14498 = n28221 & n14496 ;
  assign n14499 = n14497 | n14498 ;
  assign n14500 = n14492 & n14499 ;
  assign n15172 = n14492 | n14499 ;
  assign n31023 = ~n14500 ;
  assign n15456 = n31023 & n15172 ;
  assign n31024 = ~n15456 ;
  assign n15457 = n15455 & n31024 ;
  assign n15171 = n14511 | n15170 ;
  assign n15173 = n15171 & n15172 ;
  assign n15174 = n14500 | n15173 ;
  assign n31025 = ~n15174 ;
  assign n15458 = n15172 & n31025 ;
  assign n15459 = n15457 | n15458 ;
  assign n7214 = n3876 & n7162 ;
  assign n7157 = x[106] & n7100 ;
  assign n7725 = x[107] & n7647 ;
  assign n15460 = n7157 | n7725 ;
  assign n15461 = x[108] & n7098 ;
  assign n15462 = n15460 | n15461 ;
  assign n15463 = n7214 | n15462 ;
  assign n31026 = ~n15463 ;
  assign n15464 = x[20] & n31026 ;
  assign n15465 = n28114 & n15463 ;
  assign n15466 = n15464 | n15465 ;
  assign n31027 = ~n15466 ;
  assign n15467 = n15459 & n31027 ;
  assign n31028 = ~n15459 ;
  assign n16237 = n31028 & n15466 ;
  assign n16238 = n15467 | n16237 ;
  assign n31029 = ~n16238 ;
  assign n16347 = n16236 & n31029 ;
  assign n31030 = ~n16236 ;
  assign n16348 = n31030 & n16238 ;
  assign n16349 = n16347 | n16348 ;
  assign n8745 = n4246 & n8706 ;
  assign n8691 = x[109] & n8645 ;
  assign n9856 = x[110] & n9278 ;
  assign n16350 = n8691 | n9856 ;
  assign n16351 = x[111] & n8643 ;
  assign n16352 = n16350 | n16351 ;
  assign n16353 = n8745 | n16352 ;
  assign n31031 = ~n16353 ;
  assign n16354 = x[17] & n31031 ;
  assign n16355 = n28039 & n16353 ;
  assign n16356 = n16354 | n16355 ;
  assign n16357 = n16349 | n16356 ;
  assign n16358 = n16349 & n16356 ;
  assign n31032 = ~n16358 ;
  assign n17401 = n16357 & n31032 ;
  assign n31033 = ~n17203 ;
  assign n17402 = n31033 & n17401 ;
  assign n31034 = ~n17401 ;
  assign n17403 = n17203 & n31034 ;
  assign n17404 = n17402 | n17403 ;
  assign n17405 = n17400 & n17404 ;
  assign n18284 = n17400 | n17404 ;
  assign n31035 = ~n17405 ;
  assign n18285 = n31035 & n18284 ;
  assign n18286 = n18283 & n18285 ;
  assign n18622 = n18283 | n18285 ;
  assign n31036 = ~n18286 ;
  assign n18623 = n31036 & n18622 ;
  assign n12735 = n797 & n12695 ;
  assign n12665 = x[115] & n12633 ;
  assign n14381 = x[116] & n13533 ;
  assign n18624 = n12665 | n14381 ;
  assign n18625 = x[117] & n12631 ;
  assign n18626 = n18624 | n18625 ;
  assign n18627 = n12735 | n18626 ;
  assign n31037 = ~n18627 ;
  assign n18628 = x[11] & n31037 ;
  assign n18629 = n27892 & n18627 ;
  assign n18630 = n18628 | n18629 ;
  assign n18631 = n18623 | n18630 ;
  assign n18632 = n18623 & n18630 ;
  assign n31038 = ~n18632 ;
  assign n19907 = n18631 & n31038 ;
  assign n31039 = ~n19585 ;
  assign n19908 = n31039 & n19907 ;
  assign n31040 = ~n19907 ;
  assign n19909 = n19585 & n31040 ;
  assign n19910 = n19908 | n19909 ;
  assign n15341 = n4678 & n15308 ;
  assign n15275 = x[118] & n15246 ;
  assign n17314 = x[119] & n16288 ;
  assign n19911 = n15275 | n17314 ;
  assign n19912 = x[120] & n15244 ;
  assign n19913 = n19911 | n19912 ;
  assign n19914 = n15341 | n19913 ;
  assign n31041 = ~n19914 ;
  assign n19915 = x[8] & n31041 ;
  assign n19916 = n27845 & n19914 ;
  assign n19917 = n19915 | n19916 ;
  assign n31042 = ~n19917 ;
  assign n19918 = n19910 & n31042 ;
  assign n31043 = ~n19910 ;
  assign n19920 = n31043 & n19917 ;
  assign n19921 = n19918 | n19920 ;
  assign n18445 = n5417 & n18392 ;
  assign n18382 = x[121] & n18329 ;
  assign n18544 = x[122] & n18514 ;
  assign n19922 = n18382 | n18544 ;
  assign n19923 = x[123] & n18327 ;
  assign n19924 = n19922 | n19923 ;
  assign n19925 = n18445 | n19924 ;
  assign n31044 = ~n19925 ;
  assign n19926 = x[5] & n31044 ;
  assign n19927 = n27813 & n19925 ;
  assign n19928 = n19926 | n19927 ;
  assign n31045 = ~n19928 ;
  assign n19929 = n19921 & n31045 ;
  assign n31046 = ~n19921 ;
  assign n19951 = n31046 & n19928 ;
  assign n19952 = n19929 | n19951 ;
  assign n20928 = n19964 & n20926 ;
  assign n20929 = n19962 | n20928 ;
  assign n31047 = ~n20929 ;
  assign n20930 = n19952 & n31047 ;
  assign n31048 = ~n19952 ;
  assign n20932 = n31048 & n20929 ;
  assign n20933 = n20930 | n20932 ;
  assign n5354 = n637 & n638 ;
  assign n5355 = n27658 | n5354 ;
  assign n27273 = x[125] & x[126] ;
  assign n5356 = x[125] | x[126] ;
  assign n31049 = ~n27273 ;
  assign n5385 = n31049 & n5356 ;
  assign n5386 = n5355 & n5385 ;
  assign n5387 = n5355 | n5385 ;
  assign n31050 = ~n5386 ;
  assign n5388 = n31050 & n5387 ;
  assign n19715 = n5388 & n19656 ;
  assign n19771 = x[124] & n19723 ;
  assign n19872 = x[125] & n19829 ;
  assign n20934 = n19771 | n19872 ;
  assign n20935 = x[126] & n19655 ;
  assign n20936 = n20934 | n20935 ;
  assign n20937 = n19715 | n20936 ;
  assign n31051 = ~n20937 ;
  assign n20938 = x[2] & n31051 ;
  assign n20939 = n27790 & n20937 ;
  assign n20940 = n20938 | n20939 ;
  assign n31052 = ~n20940 ;
  assign n20941 = n20933 & n31052 ;
  assign n31053 = ~n20933 ;
  assign n20971 = n31053 & n20940 ;
  assign n20972 = n20941 | n20971 ;
  assign n20973 = n20970 & n20972 ;
  assign n23103 = n20970 | n20972 ;
  assign n31054 = ~n20973 ;
  assign n23104 = n31054 & n23103 ;
  assign n23105 = n23102 & n23104 ;
  assign n27718 = n23102 | n23104 ;
  assign n31055 = ~n23105 ;
  assign n191 = n31055 & n27718 ;
  assign n18287 = n17405 | n18286 ;
  assign n10597 = n4474 & n10542 ;
  assign n10502 = x[113] & n10481 ;
  assign n11905 = x[114] & n11232 ;
  assign n17380 = n10502 | n11905 ;
  assign n17381 = x[115] & n10479 ;
  assign n17382 = n17380 | n17381 ;
  assign n17383 = n10597 | n17382 ;
  assign n31056 = ~n17383 ;
  assign n17384 = x[14] & n31056 ;
  assign n17385 = n27956 & n17383 ;
  assign n17386 = n17384 | n17385 ;
  assign n17204 = n16357 & n17203 ;
  assign n17205 = n16358 | n17204 ;
  assign n8758 = n4442 & n8706 ;
  assign n8692 = x[110] & n8645 ;
  assign n9868 = x[111] & n9278 ;
  assign n16335 = n8692 | n9868 ;
  assign n16336 = x[112] & n8643 ;
  assign n16337 = n16335 | n16336 ;
  assign n16338 = n8758 | n16337 ;
  assign n31057 = ~n16338 ;
  assign n16339 = x[17] & n31057 ;
  assign n16340 = n28039 & n16338 ;
  assign n16341 = n16339 | n16340 ;
  assign n15468 = n15459 & n15466 ;
  assign n16239 = n16236 & n16238 ;
  assign n16240 = n15468 | n16239 ;
  assign n7193 = n3639 & n7162 ;
  assign n7144 = x[107] & n7100 ;
  assign n7724 = x[108] & n7647 ;
  assign n15437 = n7144 | n7724 ;
  assign n15438 = x[109] & n7098 ;
  assign n15439 = n15437 | n15438 ;
  assign n15440 = n7193 | n15439 ;
  assign n31058 = ~n15440 ;
  assign n15441 = x[20] & n31058 ;
  assign n15442 = n28114 & n15440 ;
  assign n15443 = n15441 | n15442 ;
  assign n5351 = n3223 & n5302 ;
  assign n5295 = x[104] & n5240 ;
  assign n6277 = x[105] & n6179 ;
  assign n14482 = n5295 | n6277 ;
  assign n14483 = x[106] & n5238 ;
  assign n14484 = n14482 | n14483 ;
  assign n14485 = n5351 | n14484 ;
  assign n31059 = ~n14485 ;
  assign n14486 = x[23] & n31059 ;
  assign n14487 = n28221 & n14485 ;
  assign n14488 = n14486 | n14487 ;
  assign n14247 = n13603 | n14246 ;
  assign n12948 = n12939 & n12946 ;
  assign n13457 = n12948 | n13456 ;
  assign n12536 = n12534 & n12535 ;
  assign n12537 = n12046 | n12536 ;
  assign n2439 = n779 & n2438 ;
  assign n686 = x[95] & n663 ;
  assign n728 = x[96] & n720 ;
  assign n12026 = n686 | n728 ;
  assign n12027 = x[97] & n652 ;
  assign n12028 = n12026 | n12027 ;
  assign n12029 = n2439 | n12028 ;
  assign n31060 = ~n12029 ;
  assign n12030 = x[32] & n31060 ;
  assign n12031 = n28658 & n12029 ;
  assign n12032 = n12030 | n12031 ;
  assign n9376 = n9367 & n9374 ;
  assign n9662 = n9376 | n9661 ;
  assign n2637 = n1239 & n2635 ;
  assign n2510 = x[83] & n2492 ;
  assign n2600 = x[84] & n2557 ;
  assign n9355 = n2510 | n2600 ;
  assign n9356 = x[85] & n2488 ;
  assign n9357 = n9355 | n9356 ;
  assign n9358 = n2637 | n9357 ;
  assign n31061 = ~n9358 ;
  assign n9359 = x[44] & n31061 ;
  assign n9360 = n29400 & n9358 ;
  assign n9361 = n9359 | n9360 ;
  assign n8882 = n8878 & n8880 ;
  assign n9114 = n9110 & n9112 ;
  assign n9115 = n8882 | n9114 ;
  assign n2010 = n1741 & n2007 ;
  assign n1923 = x[77] & n1866 ;
  assign n1982 = x[78] & n1931 ;
  assign n8267 = n1923 | n1982 ;
  assign n8268 = x[79] & n1862 ;
  assign n8269 = n8267 | n8268 ;
  assign n8270 = n2010 | n8269 ;
  assign n31062 = ~n8270 ;
  assign n8271 = x[50] & n31062 ;
  assign n8272 = n29865 & n8270 ;
  assign n8273 = n8271 | n8272 ;
  assign n7835 = n7831 & n7833 ;
  assign n7980 = n7976 & n7978 ;
  assign n7981 = n7835 | n7980 ;
  assign n7452 = n7448 & n7450 ;
  assign n7453 = n7449 | n7452 ;
  assign n3740 = n1457 & n3733 ;
  assign n1328 = x[71] & n1319 ;
  assign n1386 = x[72] & n1384 ;
  assign n7333 = n1328 | n1386 ;
  assign n7334 = x[73] & n1315 ;
  assign n7335 = n7333 | n7334 ;
  assign n7336 = n3740 | n7335 ;
  assign n31063 = ~n7336 ;
  assign n7337 = x[56] & n31063 ;
  assign n7338 = n30379 & n7336 ;
  assign n7339 = n7337 | n7338 ;
  assign n6486 = n6457 & n6484 ;
  assign n27215 = x[62] & x[63] ;
  assign n804 = x[62] | x[63] ;
  assign n31064 = ~n27215 ;
  assign n805 = n31064 & n804 ;
  assign n6487 = x[64] & n805 ;
  assign n6488 = n6486 & n6487 ;
  assign n6489 = n6486 | n6487 ;
  assign n31065 = ~n6488 ;
  assign n6490 = n31065 & n6489 ;
  assign n924 = x[65] & n900 ;
  assign n964 = x[66] & n949 ;
  assign n6491 = n924 | n964 ;
  assign n6492 = x[67] & n881 ;
  assign n6493 = n6491 | n6492 ;
  assign n6507 = n1006 & n6494 ;
  assign n6509 = n6493 | n6507 ;
  assign n31066 = ~n6509 ;
  assign n6510 = x[62] & n31066 ;
  assign n6511 = n30886 & n6509 ;
  assign n6512 = n6510 | n6511 ;
  assign n6513 = n6490 | n6512 ;
  assign n6514 = n6490 & n6512 ;
  assign n31067 = ~n6514 ;
  assign n6818 = n6513 & n31067 ;
  assign n5988 = n1217 & n5976 ;
  assign n1113 = x[68] & n1079 ;
  assign n1177 = x[69] & n1144 ;
  assign n6819 = n1113 | n1177 ;
  assign n6820 = x[70] & n1075 ;
  assign n6821 = n6819 | n6820 ;
  assign n6822 = n5988 | n6821 ;
  assign n31068 = ~n6822 ;
  assign n6823 = x[59] & n31068 ;
  assign n6824 = n30638 & n6822 ;
  assign n6825 = n6823 | n6824 ;
  assign n6826 = n6818 | n6825 ;
  assign n6827 = n6818 & n6825 ;
  assign n31069 = ~n6827 ;
  assign n6891 = n6826 & n31069 ;
  assign n6892 = n30977 & n6891 ;
  assign n31070 = ~n6891 ;
  assign n7340 = n6890 & n31070 ;
  assign n7341 = n6892 | n7340 ;
  assign n31071 = ~n7339 ;
  assign n7342 = n31071 & n7341 ;
  assign n31072 = ~n7341 ;
  assign n7454 = n7339 & n31072 ;
  assign n7455 = n7342 | n7454 ;
  assign n31073 = ~n7455 ;
  assign n7457 = n7453 & n31073 ;
  assign n31074 = ~n7453 ;
  assign n7814 = n31074 & n7455 ;
  assign n7815 = n7457 | n7814 ;
  assign n2756 = n1690 & n2750 ;
  assign n1569 = x[74] & n1551 ;
  assign n1655 = x[75] & n1616 ;
  assign n7816 = n1569 | n1655 ;
  assign n7817 = x[76] & n1547 ;
  assign n7818 = n7816 | n7817 ;
  assign n7819 = n2756 | n7818 ;
  assign n31075 = ~n7819 ;
  assign n7820 = x[53] & n31075 ;
  assign n7821 = n30125 & n7819 ;
  assign n7822 = n7820 | n7821 ;
  assign n7823 = n7815 | n7822 ;
  assign n7824 = n7815 & n7822 ;
  assign n31076 = ~n7824 ;
  assign n7982 = n7823 & n31076 ;
  assign n7983 = n7981 & n7982 ;
  assign n8274 = n7981 | n7982 ;
  assign n31077 = ~n7983 ;
  assign n8275 = n31077 & n8274 ;
  assign n8276 = n8273 & n8275 ;
  assign n8277 = n8273 | n8275 ;
  assign n31078 = ~n8276 ;
  assign n8278 = n31078 & n8277 ;
  assign n8289 = n8285 & n8287 ;
  assign n8476 = n8472 & n8474 ;
  assign n8477 = n8289 | n8476 ;
  assign n31079 = ~n8477 ;
  assign n8478 = n8278 & n31079 ;
  assign n31080 = ~n8278 ;
  assign n8861 = n31080 & n8477 ;
  assign n8862 = n8478 | n8861 ;
  assign n2342 = n1003 & n2321 ;
  assign n2238 = x[80] & n2179 ;
  assign n2269 = x[81] & n2244 ;
  assign n8863 = n2238 | n2269 ;
  assign n8864 = x[82] & n2175 ;
  assign n8865 = n8863 | n8864 ;
  assign n8866 = n2342 | n8865 ;
  assign n31081 = ~n8866 ;
  assign n8867 = x[47] & n31081 ;
  assign n8868 = n29621 & n8866 ;
  assign n8869 = n8867 | n8868 ;
  assign n8870 = n8862 | n8869 ;
  assign n8871 = n8862 & n8869 ;
  assign n31082 = ~n8871 ;
  assign n9116 = n8870 & n31082 ;
  assign n9117 = n9115 & n9116 ;
  assign n9362 = n9115 | n9116 ;
  assign n31083 = ~n9117 ;
  assign n9363 = n31083 & n9362 ;
  assign n31084 = ~n9361 ;
  assign n9364 = n31084 & n9363 ;
  assign n31085 = ~n9363 ;
  assign n9663 = n9361 & n31085 ;
  assign n9664 = n9364 | n9663 ;
  assign n9665 = n9662 & n9664 ;
  assign n10007 = n9662 | n9664 ;
  assign n31086 = ~n9665 ;
  assign n10008 = n31086 & n10007 ;
  assign n3190 = n1720 & n3162 ;
  assign n3069 = x[86] & n3031 ;
  assign n3155 = x[87] & n3096 ;
  assign n10009 = n3069 | n3155 ;
  assign n10010 = x[88] & n3027 ;
  assign n10011 = n10009 | n10010 ;
  assign n10012 = n3190 | n10011 ;
  assign n31087 = ~n10012 ;
  assign n10013 = x[41] & n31087 ;
  assign n10014 = n29184 & n10012 ;
  assign n10015 = n10013 | n10014 ;
  assign n10016 = n10008 | n10015 ;
  assign n10017 = n10008 & n10015 ;
  assign n31088 = ~n10017 ;
  assign n10018 = n10016 & n31088 ;
  assign n10354 = n10028 | n10353 ;
  assign n31089 = ~n10354 ;
  assign n10355 = n10018 & n31089 ;
  assign n31090 = ~n10018 ;
  assign n10690 = n31090 & n10354 ;
  assign n10691 = n10355 | n10690 ;
  assign n3602 = n2046 & n3574 ;
  assign n3504 = x[89] & n3443 ;
  assign n3539 = x[90] & n3508 ;
  assign n10692 = n3504 | n3539 ;
  assign n10693 = x[91] & n3439 ;
  assign n10694 = n10692 | n10693 ;
  assign n10695 = n3602 | n10694 ;
  assign n31091 = ~n10695 ;
  assign n10696 = x[38] & n31091 ;
  assign n10697 = n28996 & n10695 ;
  assign n10698 = n10696 | n10697 ;
  assign n31092 = ~n10698 ;
  assign n10699 = n10691 & n31092 ;
  assign n31093 = ~n10691 ;
  assign n10701 = n31093 & n10698 ;
  assign n10702 = n10699 | n10701 ;
  assign n10713 = n10704 & n10711 ;
  assign n11110 = n10715 & n11108 ;
  assign n11111 = n10713 | n11110 ;
  assign n31094 = ~n10702 ;
  assign n11112 = n31094 & n11111 ;
  assign n31095 = ~n11111 ;
  assign n11280 = n10702 & n31095 ;
  assign n11281 = n11112 | n11280 ;
  assign n4066 = n2410 & n4041 ;
  assign n3963 = x[92] & n3910 ;
  assign n4011 = x[93] & n3975 ;
  assign n11282 = n3963 | n4011 ;
  assign n11283 = x[94] & n3906 ;
  assign n11284 = n11282 | n11283 ;
  assign n11285 = n4066 | n11284 ;
  assign n31096 = ~n11285 ;
  assign n11286 = x[35] & n31096 ;
  assign n11287 = n28822 & n11285 ;
  assign n11288 = n11286 | n11287 ;
  assign n11289 = n11281 | n11288 ;
  assign n11290 = n11281 & n11288 ;
  assign n31097 = ~n11290 ;
  assign n11291 = n11289 & n31097 ;
  assign n11302 = n11293 & n11300 ;
  assign n11712 = n11304 & n11710 ;
  assign n11713 = n11302 | n11712 ;
  assign n11714 = n11291 & n11713 ;
  assign n12033 = n11291 | n11713 ;
  assign n31098 = ~n11714 ;
  assign n12034 = n31098 & n12033 ;
  assign n31099 = ~n12032 ;
  assign n12035 = n31099 & n12034 ;
  assign n31100 = ~n12034 ;
  assign n12538 = n12032 & n31100 ;
  assign n12539 = n12035 | n12538 ;
  assign n12540 = n12537 | n12539 ;
  assign n12541 = n12537 & n12539 ;
  assign n31101 = ~n12541 ;
  assign n12843 = n12540 & n31101 ;
  assign n4655 = n2466 & n4632 ;
  assign n4527 = x[98] & n4514 ;
  assign n4575 = x[99] & n4572 ;
  assign n12844 = n4527 | n4575 ;
  assign n12845 = x[100] & n4504 ;
  assign n12846 = n12844 | n12845 ;
  assign n12847 = n4655 | n12846 ;
  assign n31102 = ~n12847 ;
  assign n12848 = x[29] & n31102 ;
  assign n12849 = n28483 & n12847 ;
  assign n12850 = n12848 | n12849 ;
  assign n12851 = n12843 | n12850 ;
  assign n13458 = n12843 & n12850 ;
  assign n31103 = ~n13458 ;
  assign n13459 = n12851 & n31103 ;
  assign n31104 = ~n13457 ;
  assign n13460 = n31104 & n13459 ;
  assign n31105 = ~n13459 ;
  assign n13582 = n13457 & n31105 ;
  assign n13583 = n13460 | n13582 ;
  assign n2627 = n452 & n2626 ;
  assign n356 = x[101] & n330 ;
  assign n404 = x[102] & n390 ;
  assign n13584 = n356 | n404 ;
  assign n13585 = x[103] & n322 ;
  assign n13586 = n13584 | n13585 ;
  assign n13587 = n2627 | n13586 ;
  assign n31106 = ~n13587 ;
  assign n13588 = x[26] & n31106 ;
  assign n13589 = n28342 & n13587 ;
  assign n13590 = n13588 | n13589 ;
  assign n13591 = n13583 | n13590 ;
  assign n13592 = n13583 & n13590 ;
  assign n31107 = ~n13592 ;
  assign n14248 = n13591 & n31107 ;
  assign n14249 = n14247 & n14248 ;
  assign n14489 = n14247 | n14248 ;
  assign n31108 = ~n14249 ;
  assign n14490 = n31108 & n14489 ;
  assign n31109 = ~n14490 ;
  assign n15175 = n14488 & n31109 ;
  assign n31110 = ~n14488 ;
  assign n15176 = n31110 & n14490 ;
  assign n15177 = n15175 | n15176 ;
  assign n15178 = n15174 & n15177 ;
  assign n15444 = n15174 | n15176 ;
  assign n15445 = n15175 | n15444 ;
  assign n31111 = ~n15178 ;
  assign n15446 = n31111 & n15445 ;
  assign n31112 = ~n15446 ;
  assign n15447 = n15443 & n31112 ;
  assign n31113 = ~n15443 ;
  assign n16241 = n31113 & n15446 ;
  assign n16242 = n15447 | n16241 ;
  assign n16243 = n16240 & n16242 ;
  assign n16342 = n16240 | n16241 ;
  assign n16343 = n15447 | n16342 ;
  assign n31114 = ~n16243 ;
  assign n16344 = n31114 & n16343 ;
  assign n16345 = n16341 | n16344 ;
  assign n16346 = n16341 & n16344 ;
  assign n31115 = ~n16346 ;
  assign n17206 = n16345 & n31115 ;
  assign n17207 = n17205 & n17206 ;
  assign n31116 = ~n16344 ;
  assign n17387 = n16341 & n31116 ;
  assign n31117 = ~n16341 ;
  assign n17388 = n31117 & n16344 ;
  assign n17389 = n17205 | n17388 ;
  assign n17390 = n17387 | n17389 ;
  assign n31118 = ~n17207 ;
  assign n17391 = n31118 & n17390 ;
  assign n17392 = n17386 | n17391 ;
  assign n17393 = n17386 & n17391 ;
  assign n31119 = ~n17393 ;
  assign n18607 = n17392 & n31119 ;
  assign n31120 = ~n18287 ;
  assign n18608 = n31120 & n18607 ;
  assign n31121 = ~n18607 ;
  assign n18609 = n18287 & n31121 ;
  assign n18610 = n18608 | n18609 ;
  assign n12705 = n784 & n12695 ;
  assign n12669 = x[116] & n12633 ;
  assign n14393 = x[117] & n13533 ;
  assign n18611 = n12669 | n14393 ;
  assign n18612 = x[118] & n12631 ;
  assign n18613 = n18611 | n18612 ;
  assign n18614 = n12705 | n18613 ;
  assign n31122 = ~n18614 ;
  assign n18615 = x[11] & n31122 ;
  assign n18616 = n27892 & n18614 ;
  assign n18617 = n18615 | n18616 ;
  assign n31123 = ~n18617 ;
  assign n18618 = n18610 & n31123 ;
  assign n31124 = ~n18610 ;
  assign n18620 = n31124 & n18617 ;
  assign n18621 = n18618 | n18620 ;
  assign n19586 = n18631 & n19585 ;
  assign n19587 = n18632 | n19586 ;
  assign n19588 = n18621 & n19587 ;
  assign n19804 = n18621 | n19587 ;
  assign n31125 = ~n19588 ;
  assign n19805 = n31125 & n19804 ;
  assign n15346 = n4985 & n15308 ;
  assign n15277 = x[119] & n15246 ;
  assign n17316 = x[120] & n16288 ;
  assign n19806 = n15277 | n17316 ;
  assign n19807 = x[121] & n15244 ;
  assign n19808 = n19806 | n19807 ;
  assign n19809 = n15346 | n19808 ;
  assign n31126 = ~n19809 ;
  assign n19810 = x[8] & n31126 ;
  assign n19811 = n27845 & n19809 ;
  assign n19812 = n19810 | n19811 ;
  assign n19813 = n19805 | n19812 ;
  assign n19814 = n19805 & n19812 ;
  assign n31127 = ~n19814 ;
  assign n19815 = n19813 & n31127 ;
  assign n18436 = n5838 & n18392 ;
  assign n18366 = x[122] & n18329 ;
  assign n18554 = x[123] & n18514 ;
  assign n19816 = n18366 | n18554 ;
  assign n19817 = x[124] & n18327 ;
  assign n19818 = n19816 | n19817 ;
  assign n19819 = n18436 | n19818 ;
  assign n31128 = ~n19819 ;
  assign n19820 = x[5] & n31128 ;
  assign n19821 = n27813 & n19819 ;
  assign n19822 = n19820 | n19821 ;
  assign n19823 = n19815 | n19822 ;
  assign n19824 = n19815 & n19822 ;
  assign n31129 = ~n19824 ;
  assign n19906 = n19823 & n31129 ;
  assign n19919 = n19910 & n19917 ;
  assign n19930 = n19921 & n19928 ;
  assign n19931 = n19919 | n19930 ;
  assign n31130 = ~n19931 ;
  assign n19932 = n19906 & n31130 ;
  assign n31131 = ~n19906 ;
  assign n19934 = n31131 & n19931 ;
  assign n19935 = n19932 | n19934 ;
  assign n5357 = n5355 & n5356 ;
  assign n5358 = n27273 | n5357 ;
  assign n27777 = x[126] & x[127] ;
  assign n5625 = x[126] | x[127] ;
  assign n31132 = ~n27777 ;
  assign n5626 = n31132 & n5625 ;
  assign n5627 = n5358 | n5626 ;
  assign n5628 = n5358 & n5626 ;
  assign n31133 = ~n5628 ;
  assign n5629 = n5627 & n31133 ;
  assign n19671 = n5629 & n19656 ;
  assign n19768 = x[125] & n19723 ;
  assign n19873 = x[126] & n19829 ;
  assign n19936 = n19768 | n19873 ;
  assign n19937 = x[127] & n19655 ;
  assign n19938 = n19936 | n19937 ;
  assign n19939 = n19671 | n19938 ;
  assign n31134 = ~n19939 ;
  assign n19940 = x[2] & n31134 ;
  assign n19941 = n27790 & n19939 ;
  assign n19942 = n19940 | n19941 ;
  assign n31135 = ~n19942 ;
  assign n19943 = n19935 & n31135 ;
  assign n31136 = ~n19935 ;
  assign n19949 = n31136 & n19942 ;
  assign n19950 = n19943 | n19949 ;
  assign n20931 = n19952 & n20929 ;
  assign n20942 = n20933 & n20940 ;
  assign n20943 = n20931 | n20942 ;
  assign n31137 = ~n20943 ;
  assign n20944 = n19950 & n31137 ;
  assign n31138 = ~n19950 ;
  assign n20946 = n31138 & n20943 ;
  assign n20947 = n20944 | n20946 ;
  assign n23106 = n20973 | n23105 ;
  assign n23107 = n20947 | n23106 ;
  assign n23108 = n20947 & n23106 ;
  assign n31139 = ~n23108 ;
  assign n192 = n23107 & n31139 ;
  assign n20945 = n19950 & n20943 ;
  assign n23109 = n20945 | n23108 ;
  assign n19933 = n19906 & n19931 ;
  assign n19944 = n19935 & n19942 ;
  assign n19945 = n19933 | n19944 ;
  assign n31140 = ~x[127] ;
  assign n6183 = x[126] & n31140 ;
  assign n6184 = n5358 & n6183 ;
  assign n5359 = x[126] | n5358 ;
  assign n5360 = x[127] & n5359 ;
  assign n31141 = ~n5360 ;
  assign n6185 = x[127] & n31141 ;
  assign n6186 = n6184 | n6185 ;
  assign n19705 = n6186 & n19656 ;
  assign n19769 = x[126] & n19723 ;
  assign n19892 = x[127] & n19829 ;
  assign n19893 = n19769 | n19892 ;
  assign n19894 = n19705 | n19893 ;
  assign n19895 = x[2] | n19894 ;
  assign n19896 = x[2] & n19894 ;
  assign n31142 = ~n19896 ;
  assign n19897 = n19895 & n31142 ;
  assign n19825 = n19814 | n19824 ;
  assign n18619 = n18610 & n18617 ;
  assign n19589 = n18619 | n19588 ;
  assign n12727 = n5047 & n12695 ;
  assign n12677 = x[117] & n12633 ;
  assign n14363 = x[118] & n13533 ;
  assign n18597 = n12677 | n14363 ;
  assign n18598 = x[119] & n12631 ;
  assign n18599 = n18597 | n18598 ;
  assign n18600 = n12727 | n18599 ;
  assign n18601 = x[11] | n18600 ;
  assign n18602 = x[11] & n18600 ;
  assign n31143 = ~n18602 ;
  assign n18603 = n18601 & n31143 ;
  assign n18288 = n17392 & n18287 ;
  assign n18289 = n17393 | n18288 ;
  assign n10569 = n4702 & n10542 ;
  assign n10521 = x[114] & n10481 ;
  assign n11901 = x[115] & n11232 ;
  assign n17371 = n10521 | n11901 ;
  assign n17372 = x[116] & n10479 ;
  assign n17373 = n17371 | n17372 ;
  assign n17374 = n10569 | n17373 ;
  assign n17375 = x[14] | n17374 ;
  assign n17376 = x[14] & n17374 ;
  assign n31144 = ~n17376 ;
  assign n17377 = n17375 & n31144 ;
  assign n8755 = n4087 & n8706 ;
  assign n8697 = x[111] & n8645 ;
  assign n9850 = x[112] & n9278 ;
  assign n16323 = n8697 | n9850 ;
  assign n16324 = x[113] & n8643 ;
  assign n16325 = n16323 | n16324 ;
  assign n16326 = n8755 | n16325 ;
  assign n31145 = ~n16326 ;
  assign n16327 = x[17] & n31145 ;
  assign n16328 = n28039 & n16326 ;
  assign n16329 = n16327 | n16328 ;
  assign n15448 = n15443 & n15446 ;
  assign n16244 = n15448 | n16243 ;
  assign n7210 = n3615 & n7162 ;
  assign n7128 = x[108] & n7100 ;
  assign n7719 = x[109] & n7647 ;
  assign n15429 = n7128 | n7719 ;
  assign n15430 = x[110] & n7098 ;
  assign n15431 = n15429 | n15430 ;
  assign n15432 = n7210 | n15431 ;
  assign n31146 = ~n15432 ;
  assign n15433 = x[20] & n31146 ;
  assign n15434 = n28114 & n15432 ;
  assign n15435 = n15433 | n15434 ;
  assign n14491 = n14488 & n14490 ;
  assign n15179 = n14491 | n15178 ;
  assign n2842 = n779 & n2841 ;
  assign n690 = x[96] & n663 ;
  assign n730 = x[97] & n720 ;
  assign n12014 = n690 | n730 ;
  assign n12015 = x[98] & n652 ;
  assign n12016 = n12014 | n12015 ;
  assign n12017 = n2842 | n12016 ;
  assign n31147 = ~n12017 ;
  assign n12018 = x[32] & n31147 ;
  assign n12019 = n28658 & n12017 ;
  assign n12020 = n12018 | n12019 ;
  assign n2660 = n1213 & n2635 ;
  assign n2525 = x[84] & n2492 ;
  assign n2612 = x[85] & n2557 ;
  assign n9342 = n2525 | n2612 ;
  assign n9343 = x[86] & n2488 ;
  assign n9344 = n9342 | n9343 ;
  assign n9345 = n2660 | n9344 ;
  assign n31148 = ~n9345 ;
  assign n9346 = x[44] & n31148 ;
  assign n9347 = n29400 & n9345 ;
  assign n9348 = n9346 | n9347 ;
  assign n2009 = n1270 & n2007 ;
  assign n1869 = x[78] & n1866 ;
  assign n1989 = x[79] & n1931 ;
  assign n8255 = n1869 | n1989 ;
  assign n8256 = x[80] & n1862 ;
  assign n8257 = n8255 | n8256 ;
  assign n8258 = n2009 | n8257 ;
  assign n31149 = ~n8258 ;
  assign n8259 = x[50] & n31149 ;
  assign n8260 = n29865 & n8258 ;
  assign n8261 = n8259 | n8260 ;
  assign n2730 = n1457 & n2722 ;
  assign n1353 = x[72] & n1319 ;
  assign n1441 = x[73] & n1384 ;
  assign n7320 = n1353 | n1441 ;
  assign n7321 = x[74] & n1315 ;
  assign n7322 = n7320 | n7321 ;
  assign n7323 = n2730 | n7322 ;
  assign n31150 = ~n7323 ;
  assign n7324 = x[56] & n31150 ;
  assign n7325 = n30379 & n7323 ;
  assign n7326 = n7324 | n7325 ;
  assign n6893 = n6890 & n6891 ;
  assign n6894 = n6827 | n6893 ;
  assign n6401 = x[65] & n805 ;
  assign n6402 = x[64] & n27215 ;
  assign n6403 = n6401 | n6402 ;
  assign n908 = x[66] & n900 ;
  assign n951 = x[67] & n949 ;
  assign n6404 = n908 | n951 ;
  assign n6405 = x[68] & n881 ;
  assign n6406 = n6404 | n6405 ;
  assign n6413 = n1006 & n6408 ;
  assign n6423 = n6406 | n6413 ;
  assign n31151 = ~n6423 ;
  assign n6424 = x[62] & n31151 ;
  assign n6425 = n30886 & n6423 ;
  assign n6426 = n6424 | n6425 ;
  assign n31152 = ~n6426 ;
  assign n6427 = n6403 & n31152 ;
  assign n31153 = ~n6403 ;
  assign n6429 = n31153 & n6426 ;
  assign n6430 = n6427 | n6429 ;
  assign n6515 = n6488 | n6514 ;
  assign n31154 = ~n6515 ;
  assign n6516 = n6430 & n31154 ;
  assign n31155 = ~n6430 ;
  assign n6807 = n31155 & n6515 ;
  assign n6808 = n6516 | n6807 ;
  assign n4803 = n1217 & n4790 ;
  assign n1138 = x[69] & n1079 ;
  assign n1197 = x[70] & n1144 ;
  assign n6809 = n1138 | n1197 ;
  assign n6810 = x[71] & n1075 ;
  assign n6811 = n6809 | n6810 ;
  assign n6812 = n4803 | n6811 ;
  assign n31156 = ~n6812 ;
  assign n6813 = x[59] & n31156 ;
  assign n6814 = n30638 & n6812 ;
  assign n6815 = n6813 | n6814 ;
  assign n31157 = ~n6815 ;
  assign n6816 = n6808 & n31157 ;
  assign n31158 = ~n6808 ;
  assign n6895 = n31158 & n6815 ;
  assign n6896 = n6816 | n6895 ;
  assign n31159 = ~n6894 ;
  assign n6897 = n31159 & n6896 ;
  assign n31160 = ~n6896 ;
  assign n7327 = n6894 & n31160 ;
  assign n7328 = n6897 | n7327 ;
  assign n31161 = ~n7326 ;
  assign n7329 = n31161 & n7328 ;
  assign n31162 = ~n7328 ;
  assign n7331 = n7326 & n31162 ;
  assign n7332 = n7329 | n7331 ;
  assign n7343 = n7339 & n7341 ;
  assign n7456 = n7453 & n7455 ;
  assign n7458 = n7343 | n7456 ;
  assign n7459 = n7332 | n7458 ;
  assign n7460 = n7332 & n7458 ;
  assign n31163 = ~n7460 ;
  assign n7802 = n7459 & n31163 ;
  assign n1778 = n1690 & n1775 ;
  assign n1591 = x[75] & n1551 ;
  assign n1647 = x[76] & n1616 ;
  assign n7803 = n1591 | n1647 ;
  assign n7804 = x[77] & n1547 ;
  assign n7805 = n7803 | n7804 ;
  assign n7806 = n1778 | n7805 ;
  assign n31164 = ~n7806 ;
  assign n7807 = x[53] & n31164 ;
  assign n7808 = n30125 & n7806 ;
  assign n7809 = n7807 | n7808 ;
  assign n31165 = ~n7809 ;
  assign n7810 = n7802 & n31165 ;
  assign n31166 = ~n7802 ;
  assign n7812 = n31166 & n7809 ;
  assign n7813 = n7810 | n7812 ;
  assign n7984 = n7824 | n7983 ;
  assign n7985 = n7813 | n7984 ;
  assign n7986 = n7813 & n7984 ;
  assign n31167 = ~n7986 ;
  assign n8262 = n7985 & n31167 ;
  assign n31168 = ~n8261 ;
  assign n8263 = n31168 & n8262 ;
  assign n31169 = ~n8262 ;
  assign n8265 = n8261 & n31169 ;
  assign n8266 = n8263 | n8265 ;
  assign n8479 = n8278 & n8477 ;
  assign n8480 = n8276 | n8479 ;
  assign n8481 = n8266 | n8480 ;
  assign n8482 = n8266 & n8480 ;
  assign n31170 = ~n8482 ;
  assign n8849 = n8481 & n31170 ;
  assign n2324 = n1057 & n2321 ;
  assign n2210 = x[81] & n2179 ;
  assign n2302 = x[82] & n2244 ;
  assign n8850 = n2210 | n2302 ;
  assign n8851 = x[83] & n2175 ;
  assign n8852 = n8850 | n8851 ;
  assign n8853 = n2324 | n8852 ;
  assign n31171 = ~n8853 ;
  assign n8854 = x[47] & n31171 ;
  assign n8855 = n29621 & n8853 ;
  assign n8856 = n8854 | n8855 ;
  assign n31172 = ~n8856 ;
  assign n8857 = n8849 & n31172 ;
  assign n31173 = ~n8849 ;
  assign n8859 = n31173 & n8856 ;
  assign n8860 = n8857 | n8859 ;
  assign n9118 = n8871 | n9117 ;
  assign n31174 = ~n9118 ;
  assign n9119 = n8860 & n31174 ;
  assign n31175 = ~n8860 ;
  assign n9349 = n31175 & n9118 ;
  assign n9350 = n9119 | n9349 ;
  assign n31176 = ~n9348 ;
  assign n9351 = n31176 & n9350 ;
  assign n31177 = ~n9350 ;
  assign n9353 = n9348 & n31177 ;
  assign n9354 = n9351 | n9353 ;
  assign n9365 = n9361 & n9363 ;
  assign n9666 = n9365 | n9665 ;
  assign n31178 = ~n9666 ;
  assign n9667 = n9354 & n31178 ;
  assign n31179 = ~n9354 ;
  assign n9995 = n31179 & n9666 ;
  assign n9996 = n9667 | n9995 ;
  assign n3171 = n1453 & n3162 ;
  assign n3062 = x[87] & n3031 ;
  assign n3139 = x[88] & n3096 ;
  assign n9997 = n3062 | n3139 ;
  assign n9998 = x[89] & n3027 ;
  assign n9999 = n9997 | n9998 ;
  assign n10000 = n3171 | n9999 ;
  assign n31180 = ~n10000 ;
  assign n10001 = x[41] & n31180 ;
  assign n10002 = n29184 & n10000 ;
  assign n10003 = n10001 | n10002 ;
  assign n10004 = n9996 | n10003 ;
  assign n10005 = n9996 & n10003 ;
  assign n31181 = ~n10005 ;
  assign n10006 = n10004 & n31181 ;
  assign n10356 = n10018 & n10354 ;
  assign n10357 = n10017 | n10356 ;
  assign n31182 = ~n10357 ;
  assign n10358 = n10006 & n31182 ;
  assign n31183 = ~n10006 ;
  assign n10677 = n31183 & n10357 ;
  assign n10678 = n10358 | n10677 ;
  assign n3610 = n1841 & n3574 ;
  assign n3502 = x[90] & n3443 ;
  assign n3558 = x[91] & n3508 ;
  assign n10679 = n3502 | n3558 ;
  assign n10680 = x[92] & n3439 ;
  assign n10681 = n10679 | n10680 ;
  assign n10682 = n3610 | n10681 ;
  assign n31184 = ~n10682 ;
  assign n10683 = x[38] & n31184 ;
  assign n10684 = n28996 & n10682 ;
  assign n10685 = n10683 | n10684 ;
  assign n31185 = ~n10685 ;
  assign n10686 = n10678 & n31185 ;
  assign n31186 = ~n10678 ;
  assign n10688 = n31186 & n10685 ;
  assign n10689 = n10686 | n10688 ;
  assign n10700 = n10691 & n10698 ;
  assign n11113 = n10702 & n11111 ;
  assign n11114 = n10700 | n11113 ;
  assign n31187 = ~n10689 ;
  assign n11115 = n31187 & n11114 ;
  assign n31188 = ~n11114 ;
  assign n11268 = n10689 & n31188 ;
  assign n11269 = n11115 | n11268 ;
  assign n4076 = n2152 & n4041 ;
  assign n3960 = x[93] & n3910 ;
  assign n4025 = x[94] & n3975 ;
  assign n11270 = n3960 | n4025 ;
  assign n11271 = x[95] & n3906 ;
  assign n11272 = n11270 | n11271 ;
  assign n11273 = n4076 | n11272 ;
  assign n31189 = ~n11273 ;
  assign n11274 = x[35] & n31189 ;
  assign n11275 = n28822 & n11273 ;
  assign n11276 = n11274 | n11275 ;
  assign n11277 = n11269 | n11276 ;
  assign n11278 = n11269 & n11276 ;
  assign n31190 = ~n11278 ;
  assign n11279 = n11277 & n31190 ;
  assign n11715 = n11290 | n11714 ;
  assign n31191 = ~n11715 ;
  assign n11716 = n11279 & n31191 ;
  assign n31192 = ~n11279 ;
  assign n12021 = n31192 & n11715 ;
  assign n12022 = n11716 | n12021 ;
  assign n12023 = n12020 | n12022 ;
  assign n12024 = n12020 & n12022 ;
  assign n31193 = ~n12024 ;
  assign n12025 = n12023 & n31193 ;
  assign n12036 = n12032 & n12034 ;
  assign n12542 = n12036 | n12541 ;
  assign n31194 = ~n12542 ;
  assign n12543 = n12025 & n31194 ;
  assign n31195 = ~n12025 ;
  assign n12831 = n31195 & n12542 ;
  assign n12832 = n12543 | n12831 ;
  assign n4643 = n2977 & n4632 ;
  assign n4534 = x[99] & n4514 ;
  assign n4584 = x[100] & n4572 ;
  assign n12833 = n4534 | n4584 ;
  assign n12834 = x[101] & n4504 ;
  assign n12835 = n12833 | n12834 ;
  assign n12836 = n4643 | n12835 ;
  assign n31196 = ~n12836 ;
  assign n12837 = x[29] & n31196 ;
  assign n12838 = n28483 & n12836 ;
  assign n12839 = n12837 | n12838 ;
  assign n12840 = n12832 | n12839 ;
  assign n12841 = n12832 & n12839 ;
  assign n31197 = ~n12841 ;
  assign n12842 = n12840 & n31197 ;
  assign n13461 = n13457 & n13459 ;
  assign n13462 = n13458 | n13461 ;
  assign n13463 = n12842 & n13462 ;
  assign n13570 = n12842 | n13462 ;
  assign n31198 = ~n13463 ;
  assign n13571 = n31198 & n13570 ;
  assign n3004 = n452 & n3001 ;
  assign n383 = x[102] & n330 ;
  assign n422 = x[103] & n390 ;
  assign n13572 = n383 | n422 ;
  assign n13573 = x[104] & n322 ;
  assign n13574 = n13572 | n13573 ;
  assign n13575 = n3004 | n13574 ;
  assign n31199 = ~n13575 ;
  assign n13576 = x[26] & n31199 ;
  assign n13577 = n28342 & n13575 ;
  assign n13578 = n13576 | n13577 ;
  assign n13579 = n13571 | n13578 ;
  assign n13580 = n13571 & n13578 ;
  assign n31200 = ~n13580 ;
  assign n13581 = n13579 & n31200 ;
  assign n14250 = n13592 | n14249 ;
  assign n31201 = ~n14250 ;
  assign n14251 = n13581 & n31201 ;
  assign n31202 = ~n13581 ;
  assign n15180 = n31202 & n14250 ;
  assign n15181 = n14251 | n15180 ;
  assign n5353 = n3199 & n5302 ;
  assign n5301 = x[105] & n5240 ;
  assign n6281 = x[106] & n6179 ;
  assign n15182 = n5301 | n6281 ;
  assign n15183 = x[107] & n5238 ;
  assign n15184 = n15182 | n15183 ;
  assign n15185 = n5353 | n15184 ;
  assign n31203 = ~n15185 ;
  assign n15186 = x[23] & n31203 ;
  assign n15187 = n28221 & n15185 ;
  assign n15188 = n15186 | n15187 ;
  assign n15189 = n15181 | n15188 ;
  assign n15190 = n15181 & n15188 ;
  assign n31204 = ~n15190 ;
  assign n15191 = n15189 & n31204 ;
  assign n15192 = n15179 | n15191 ;
  assign n15193 = n15179 & n15191 ;
  assign n31205 = ~n15193 ;
  assign n15436 = n15192 & n31205 ;
  assign n31206 = ~n15436 ;
  assign n16245 = n15435 & n31206 ;
  assign n31207 = ~n15435 ;
  assign n16246 = n31207 & n15436 ;
  assign n16247 = n16245 | n16246 ;
  assign n16248 = n16244 & n16247 ;
  assign n16330 = n16244 | n16246 ;
  assign n16331 = n16245 | n16330 ;
  assign n31208 = ~n16248 ;
  assign n16332 = n31208 & n16331 ;
  assign n31209 = ~n16332 ;
  assign n16333 = n16329 & n31209 ;
  assign n17208 = n16346 | n17207 ;
  assign n31210 = ~n16329 ;
  assign n17209 = n31210 & n16332 ;
  assign n17210 = n17208 | n17209 ;
  assign n17211 = n16333 | n17210 ;
  assign n17212 = n16333 | n17209 ;
  assign n17213 = n17208 & n17212 ;
  assign n31211 = ~n17213 ;
  assign n17378 = n17211 & n31211 ;
  assign n17379 = n17377 & n17378 ;
  assign n18290 = n17377 | n17378 ;
  assign n31212 = ~n17379 ;
  assign n18291 = n31212 & n18290 ;
  assign n31213 = ~n18291 ;
  assign n18292 = n18289 & n31213 ;
  assign n31214 = ~n18289 ;
  assign n18604 = n31214 & n18291 ;
  assign n18605 = n18292 | n18604 ;
  assign n18606 = n18603 & n18605 ;
  assign n19590 = n18603 | n18605 ;
  assign n31215 = ~n18606 ;
  assign n19591 = n31215 & n19590 ;
  assign n31216 = ~n19589 ;
  assign n19592 = n31216 & n19591 ;
  assign n31217 = ~n19591 ;
  assign n19630 = n19589 & n31217 ;
  assign n19631 = n19592 | n19630 ;
  assign n15347 = n5022 & n15308 ;
  assign n15263 = x[120] & n15246 ;
  assign n17315 = x[121] & n16288 ;
  assign n19632 = n15263 | n17315 ;
  assign n19633 = x[122] & n15244 ;
  assign n19634 = n19632 | n19633 ;
  assign n19635 = n15347 | n19634 ;
  assign n31218 = ~n19635 ;
  assign n19636 = x[8] & n31218 ;
  assign n19637 = n27845 & n19635 ;
  assign n19638 = n19636 | n19637 ;
  assign n31219 = ~n19638 ;
  assign n19639 = n19631 & n31219 ;
  assign n31220 = ~n19631 ;
  assign n19641 = n31220 & n19638 ;
  assign n19642 = n19639 | n19641 ;
  assign n18438 = n642 & n18392 ;
  assign n18348 = x[123] & n18329 ;
  assign n18549 = x[124] & n18514 ;
  assign n19643 = n18348 | n18549 ;
  assign n19644 = x[125] & n18327 ;
  assign n19645 = n19643 | n19644 ;
  assign n19646 = n18438 | n19645 ;
  assign n31221 = ~n19646 ;
  assign n19647 = x[5] & n31221 ;
  assign n19648 = n27813 & n19646 ;
  assign n19649 = n19647 | n19648 ;
  assign n19650 = n19642 | n19649 ;
  assign n19651 = n19642 & n19649 ;
  assign n31222 = ~n19651 ;
  assign n19826 = n19650 & n31222 ;
  assign n31223 = ~n19826 ;
  assign n19827 = n19825 & n31223 ;
  assign n31224 = ~n19825 ;
  assign n19898 = n31224 & n19826 ;
  assign n19899 = n19827 | n19898 ;
  assign n19900 = n19897 & n19899 ;
  assign n19946 = n19897 | n19899 ;
  assign n31225 = ~n19900 ;
  assign n19947 = n31225 & n19946 ;
  assign n19948 = n19945 & n19947 ;
  assign n23110 = n19945 | n19947 ;
  assign n31226 = ~n19948 ;
  assign n23111 = n31226 & n23110 ;
  assign n23112 = n23109 & n23111 ;
  assign n27721 = n23109 | n23111 ;
  assign n31227 = ~n23112 ;
  assign n193 = n31227 & n27721 ;
  assign n10588 = n797 & n10542 ;
  assign n10527 = x[115] & n10481 ;
  assign n11895 = x[116] & n11232 ;
  assign n17359 = n10527 | n11895 ;
  assign n17360 = x[117] & n10479 ;
  assign n17361 = n17359 | n17360 ;
  assign n17362 = n10588 | n17361 ;
  assign n17363 = x[14] | n17362 ;
  assign n17364 = x[14] & n17362 ;
  assign n31228 = ~n17364 ;
  assign n17365 = n17363 & n31228 ;
  assign n16334 = n16329 & n16332 ;
  assign n17214 = n16334 | n17213 ;
  assign n16249 = n15435 & n15436 ;
  assign n16250 = n16248 | n16249 ;
  assign n7213 = n4246 & n7162 ;
  assign n7151 = x[109] & n7100 ;
  assign n7715 = x[110] & n7647 ;
  assign n15418 = n7151 | n7715 ;
  assign n15419 = x[111] & n7098 ;
  assign n15420 = n15418 | n15419 ;
  assign n15421 = n7213 | n15420 ;
  assign n31229 = ~n15421 ;
  assign n15422 = x[20] & n31229 ;
  assign n15423 = n28114 & n15421 ;
  assign n15424 = n15422 | n15423 ;
  assign n14252 = n13581 & n14250 ;
  assign n14253 = n13580 | n14252 ;
  assign n9352 = n9348 & n9350 ;
  assign n9668 = n9354 & n9666 ;
  assign n9669 = n9352 | n9668 ;
  assign n8858 = n8849 & n8856 ;
  assign n9120 = n8860 & n9118 ;
  assign n9121 = n8858 | n9120 ;
  assign n8264 = n8261 & n8262 ;
  assign n8483 = n8264 | n8482 ;
  assign n7811 = n7802 & n7809 ;
  assign n7987 = n7811 | n7986 ;
  assign n2088 = n1690 & n2084 ;
  assign n1603 = x[76] & n1551 ;
  assign n1645 = x[77] & n1616 ;
  assign n7792 = n1603 | n1645 ;
  assign n7793 = x[78] & n1547 ;
  assign n7794 = n7792 | n7793 ;
  assign n7795 = n2088 | n7794 ;
  assign n7796 = x[53] | n7795 ;
  assign n7797 = x[53] & n7795 ;
  assign n31230 = ~n7797 ;
  assign n7798 = n7796 & n31230 ;
  assign n7330 = n7326 & n7328 ;
  assign n7461 = n7330 | n7460 ;
  assign n6817 = n6808 & n6815 ;
  assign n6898 = n6894 & n6896 ;
  assign n6899 = n6817 | n6898 ;
  assign n257 = x[65] & n27215 ;
  assign n852 = x[66] & n805 ;
  assign n6375 = n257 | n852 ;
  assign n909 = x[67] & n900 ;
  assign n977 = x[68] & n949 ;
  assign n6376 = n909 | n977 ;
  assign n6377 = x[69] & n881 ;
  assign n6378 = n6376 | n6377 ;
  assign n6392 = n1006 & n6379 ;
  assign n6394 = n6378 | n6392 ;
  assign n31231 = ~n6394 ;
  assign n6395 = x[62] & n31231 ;
  assign n6396 = n30886 & n6394 ;
  assign n6397 = n6395 | n6396 ;
  assign n6398 = n6375 | n6397 ;
  assign n6399 = n6375 & n6397 ;
  assign n31232 = ~n6399 ;
  assign n6400 = n6398 & n31232 ;
  assign n6428 = n6403 & n6426 ;
  assign n6517 = n6430 & n6515 ;
  assign n6518 = n6428 | n6517 ;
  assign n6519 = n6400 | n6518 ;
  assign n6520 = n6400 & n6518 ;
  assign n31233 = ~n6520 ;
  assign n6798 = n6519 & n31233 ;
  assign n3711 = n1217 & n3701 ;
  assign n1082 = x[70] & n1079 ;
  assign n1202 = x[71] & n1144 ;
  assign n6799 = n1082 | n1202 ;
  assign n6800 = x[72] & n1075 ;
  assign n6801 = n6799 | n6800 ;
  assign n6802 = n3711 | n6801 ;
  assign n31234 = ~n6802 ;
  assign n6803 = x[59] & n31234 ;
  assign n6804 = n30638 & n6802 ;
  assign n6805 = n6803 | n6804 ;
  assign n6806 = n6798 & n6805 ;
  assign n6900 = n6798 | n6805 ;
  assign n31235 = ~n6806 ;
  assign n6901 = n31235 & n6900 ;
  assign n31236 = ~n6901 ;
  assign n7309 = n6899 & n31236 ;
  assign n6902 = n6899 & n6900 ;
  assign n6903 = n6806 | n6902 ;
  assign n31237 = ~n6903 ;
  assign n7310 = n6900 & n31237 ;
  assign n7311 = n7309 | n7310 ;
  assign n3297 = n1457 & n3289 ;
  assign n1356 = x[73] & n1319 ;
  assign n1430 = x[74] & n1384 ;
  assign n7312 = n1356 | n1430 ;
  assign n7313 = x[75] & n1315 ;
  assign n7314 = n7312 | n7313 ;
  assign n7315 = n3297 | n7314 ;
  assign n31238 = ~n7315 ;
  assign n7316 = x[56] & n31238 ;
  assign n7317 = n30379 & n7315 ;
  assign n7318 = n7316 | n7317 ;
  assign n7319 = n7311 | n7318 ;
  assign n7462 = n7311 & n7318 ;
  assign n31239 = ~n7462 ;
  assign n7463 = n7319 & n31239 ;
  assign n31240 = ~n7461 ;
  assign n7464 = n31240 & n7463 ;
  assign n31241 = ~n7463 ;
  assign n7799 = n7461 & n31241 ;
  assign n7800 = n7464 | n7799 ;
  assign n7801 = n7798 & n7800 ;
  assign n7988 = n7798 | n7800 ;
  assign n31242 = ~n7801 ;
  assign n7989 = n31242 & n7988 ;
  assign n31243 = ~n7989 ;
  assign n7990 = n7987 & n31243 ;
  assign n31244 = ~n7987 ;
  assign n8244 = n31244 & n7989 ;
  assign n8245 = n7990 | n8244 ;
  assign n2013 = n1029 & n2007 ;
  assign n1920 = x[79] & n1866 ;
  assign n1976 = x[80] & n1931 ;
  assign n8246 = n1920 | n1976 ;
  assign n8247 = x[81] & n1862 ;
  assign n8248 = n8246 | n8247 ;
  assign n8249 = n2013 | n8248 ;
  assign n31245 = ~n8249 ;
  assign n8250 = x[50] & n31245 ;
  assign n8251 = n29865 & n8249 ;
  assign n8252 = n8250 | n8251 ;
  assign n8253 = n8245 | n8252 ;
  assign n8254 = n8245 & n8252 ;
  assign n31246 = ~n8254 ;
  assign n8484 = n8253 & n31246 ;
  assign n8485 = n8483 & n8484 ;
  assign n8838 = n8483 | n8484 ;
  assign n31247 = ~n8485 ;
  assign n8839 = n31247 & n8838 ;
  assign n2333 = n1293 & n2321 ;
  assign n2225 = x[82] & n2179 ;
  assign n2300 = x[83] & n2244 ;
  assign n8840 = n2225 | n2300 ;
  assign n8841 = x[84] & n2175 ;
  assign n8842 = n8840 | n8841 ;
  assign n8843 = n2333 | n8842 ;
  assign n31248 = ~n8843 ;
  assign n8844 = x[47] & n31248 ;
  assign n8845 = n29621 & n8843 ;
  assign n8846 = n8844 | n8845 ;
  assign n31249 = ~n8846 ;
  assign n8847 = n8839 & n31249 ;
  assign n31250 = ~n8839 ;
  assign n9122 = n31250 & n8846 ;
  assign n9123 = n8847 | n9122 ;
  assign n31251 = ~n9123 ;
  assign n9125 = n9121 & n31251 ;
  assign n31252 = ~n9121 ;
  assign n9331 = n31252 & n9123 ;
  assign n9332 = n9125 | n9331 ;
  assign n2659 = n1522 & n2635 ;
  assign n2551 = x[85] & n2492 ;
  assign n2611 = x[86] & n2557 ;
  assign n9333 = n2551 | n2611 ;
  assign n9334 = x[87] & n2488 ;
  assign n9335 = n9333 | n9334 ;
  assign n9336 = n2659 | n9335 ;
  assign n31253 = ~n9336 ;
  assign n9337 = x[44] & n31253 ;
  assign n9338 = n29400 & n9336 ;
  assign n9339 = n9337 | n9338 ;
  assign n9340 = n9332 | n9339 ;
  assign n9341 = n9332 & n9339 ;
  assign n31254 = ~n9341 ;
  assign n9670 = n9340 & n31254 ;
  assign n9671 = n9669 & n9670 ;
  assign n9982 = n9669 | n9670 ;
  assign n31255 = ~n9671 ;
  assign n9983 = n31255 & n9982 ;
  assign n3165 = n1482 & n3162 ;
  assign n3081 = x[88] & n3031 ;
  assign n3126 = x[89] & n3096 ;
  assign n9984 = n3081 | n3126 ;
  assign n9985 = x[90] & n3027 ;
  assign n9986 = n9984 | n9985 ;
  assign n9987 = n3165 | n9986 ;
  assign n31256 = ~n9987 ;
  assign n9988 = x[41] & n31256 ;
  assign n9989 = n29184 & n9987 ;
  assign n9990 = n9988 | n9989 ;
  assign n31257 = ~n9990 ;
  assign n9991 = n9983 & n31257 ;
  assign n31258 = ~n9983 ;
  assign n9993 = n31258 & n9990 ;
  assign n9994 = n9991 | n9993 ;
  assign n10359 = n10006 & n10357 ;
  assign n10360 = n10005 | n10359 ;
  assign n31259 = ~n10360 ;
  assign n10361 = n9994 & n31259 ;
  assign n31260 = ~n9994 ;
  assign n10664 = n31260 & n10360 ;
  assign n10665 = n10361 | n10664 ;
  assign n3584 = n1685 & n3574 ;
  assign n3485 = x[91] & n3443 ;
  assign n3568 = x[92] & n3508 ;
  assign n10666 = n3485 | n3568 ;
  assign n10667 = x[93] & n3439 ;
  assign n10668 = n10666 | n10667 ;
  assign n10669 = n3584 | n10668 ;
  assign n31261 = ~n10669 ;
  assign n10670 = x[38] & n31261 ;
  assign n10671 = n28996 & n10669 ;
  assign n10672 = n10670 | n10671 ;
  assign n31262 = ~n10672 ;
  assign n10673 = n10665 & n31262 ;
  assign n31263 = ~n10665 ;
  assign n10675 = n31263 & n10672 ;
  assign n10676 = n10673 | n10675 ;
  assign n10687 = n10678 & n10685 ;
  assign n11116 = n10689 & n11114 ;
  assign n11117 = n10687 | n11116 ;
  assign n31264 = ~n11117 ;
  assign n11118 = n10676 & n31264 ;
  assign n31265 = ~n10676 ;
  assign n11258 = n31265 & n11117 ;
  assign n11259 = n11118 | n11258 ;
  assign n4075 = n2000 & n4041 ;
  assign n3961 = x[94] & n3910 ;
  assign n4006 = x[95] & n3975 ;
  assign n11260 = n3961 | n4006 ;
  assign n11261 = x[96] & n3906 ;
  assign n11262 = n11260 | n11261 ;
  assign n11263 = n4075 | n11262 ;
  assign n31266 = ~n11263 ;
  assign n11264 = x[35] & n31266 ;
  assign n11265 = n28822 & n11263 ;
  assign n11266 = n11264 | n11265 ;
  assign n11719 = n11259 | n11266 ;
  assign n11267 = n11259 & n11266 ;
  assign n11717 = n11279 & n11715 ;
  assign n11718 = n11278 | n11717 ;
  assign n11720 = n11718 & n11719 ;
  assign n11721 = n11267 | n11720 ;
  assign n31267 = ~n11721 ;
  assign n11722 = n11719 & n31267 ;
  assign n31268 = ~n11267 ;
  assign n12001 = n31268 & n11719 ;
  assign n31269 = ~n12001 ;
  assign n12002 = n11718 & n31269 ;
  assign n12003 = n11722 | n12002 ;
  assign n2318 = n779 & n2313 ;
  assign n675 = x[97] & n663 ;
  assign n732 = x[98] & n720 ;
  assign n12004 = n675 | n732 ;
  assign n12005 = x[99] & n652 ;
  assign n12006 = n12004 | n12005 ;
  assign n12007 = n2318 | n12006 ;
  assign n31270 = ~n12007 ;
  assign n12008 = x[32] & n31270 ;
  assign n12009 = n28658 & n12007 ;
  assign n12010 = n12008 | n12009 ;
  assign n12011 = n12003 | n12010 ;
  assign n12012 = n12003 & n12010 ;
  assign n31271 = ~n12012 ;
  assign n12013 = n12011 & n31271 ;
  assign n12544 = n12025 & n12542 ;
  assign n12545 = n12024 | n12544 ;
  assign n12546 = n12013 | n12545 ;
  assign n12547 = n12013 & n12545 ;
  assign n31272 = ~n12547 ;
  assign n12819 = n12546 & n31272 ;
  assign n4663 = n2867 & n4632 ;
  assign n4520 = x[100] & n4514 ;
  assign n4599 = x[101] & n4572 ;
  assign n12820 = n4520 | n4599 ;
  assign n12821 = x[102] & n4504 ;
  assign n12822 = n12820 | n12821 ;
  assign n12823 = n4663 | n12822 ;
  assign n31273 = ~n12823 ;
  assign n12824 = x[29] & n31273 ;
  assign n12825 = n28483 & n12823 ;
  assign n12826 = n12824 | n12825 ;
  assign n31274 = ~n12826 ;
  assign n12827 = n12819 & n31274 ;
  assign n31275 = ~n12819 ;
  assign n12829 = n31275 & n12826 ;
  assign n12830 = n12827 | n12829 ;
  assign n13464 = n12841 | n13463 ;
  assign n31276 = ~n13464 ;
  assign n13465 = n12830 & n31276 ;
  assign n31277 = ~n12830 ;
  assign n13560 = n31277 & n13464 ;
  assign n13561 = n13465 | n13560 ;
  assign n3414 = n452 & n3409 ;
  assign n364 = x[103] & n330 ;
  assign n398 = x[104] & n390 ;
  assign n13562 = n364 | n398 ;
  assign n13563 = x[105] & n322 ;
  assign n13564 = n13562 | n13563 ;
  assign n13565 = n3414 | n13564 ;
  assign n31278 = ~n13565 ;
  assign n13566 = x[26] & n31278 ;
  assign n13567 = n28342 & n13565 ;
  assign n13568 = n13566 | n13567 ;
  assign n13569 = n13561 & n13568 ;
  assign n14254 = n13561 | n13568 ;
  assign n31279 = ~n13569 ;
  assign n14467 = n31279 & n14254 ;
  assign n31280 = ~n14467 ;
  assign n14468 = n14253 & n31280 ;
  assign n14255 = n14253 & n14254 ;
  assign n14256 = n13569 | n14255 ;
  assign n31281 = ~n14256 ;
  assign n14469 = n14254 & n31281 ;
  assign n14470 = n14468 | n14469 ;
  assign n5350 = n3876 & n5302 ;
  assign n5292 = x[106] & n5240 ;
  assign n6267 = x[107] & n6179 ;
  assign n14471 = n5292 | n6267 ;
  assign n14472 = x[108] & n5238 ;
  assign n14473 = n14471 | n14472 ;
  assign n14474 = n5350 | n14473 ;
  assign n31282 = ~n14474 ;
  assign n14475 = x[23] & n31282 ;
  assign n14476 = n28221 & n14474 ;
  assign n14477 = n14475 | n14476 ;
  assign n31283 = ~n14477 ;
  assign n14478 = n14470 & n31283 ;
  assign n31284 = ~n14470 ;
  assign n14480 = n31284 & n14477 ;
  assign n14481 = n14478 | n14480 ;
  assign n15194 = n15190 | n15193 ;
  assign n31285 = ~n15194 ;
  assign n15195 = n14481 & n31285 ;
  assign n31286 = ~n14481 ;
  assign n15425 = n31286 & n15194 ;
  assign n15426 = n15195 | n15425 ;
  assign n31287 = ~n15424 ;
  assign n15427 = n31287 & n15426 ;
  assign n31288 = ~n15426 ;
  assign n16251 = n15424 & n31288 ;
  assign n16252 = n15427 | n16251 ;
  assign n31289 = ~n16252 ;
  assign n16253 = n16250 & n31289 ;
  assign n31290 = ~n16250 ;
  assign n16313 = n31290 & n16252 ;
  assign n16314 = n16253 | n16313 ;
  assign n8752 = n4276 & n8706 ;
  assign n8677 = x[112] & n8645 ;
  assign n9877 = x[113] & n9278 ;
  assign n16315 = n8677 | n9877 ;
  assign n16316 = x[114] & n8643 ;
  assign n16317 = n16315 | n16316 ;
  assign n16318 = n8752 | n16317 ;
  assign n31291 = ~n16318 ;
  assign n16319 = x[17] & n31291 ;
  assign n16320 = n28039 & n16318 ;
  assign n16321 = n16319 | n16320 ;
  assign n16322 = n16314 | n16321 ;
  assign n17215 = n16314 & n16321 ;
  assign n31292 = ~n17215 ;
  assign n17216 = n16322 & n31292 ;
  assign n17217 = n17214 & n17216 ;
  assign n17366 = n17214 | n17216 ;
  assign n31293 = ~n17217 ;
  assign n17367 = n31293 & n17366 ;
  assign n17368 = n17365 & n17367 ;
  assign n17369 = n17365 | n17367 ;
  assign n31294 = ~n17368 ;
  assign n17370 = n31294 & n17369 ;
  assign n18293 = n18289 & n18291 ;
  assign n18294 = n17379 | n18293 ;
  assign n18295 = n17370 & n18294 ;
  assign n18484 = n17370 | n18294 ;
  assign n31295 = ~n18295 ;
  assign n18485 = n31295 & n18484 ;
  assign n12724 = n4678 & n12695 ;
  assign n12670 = x[118] & n12633 ;
  assign n14398 = x[119] & n13533 ;
  assign n18486 = n12670 | n14398 ;
  assign n18487 = x[120] & n12631 ;
  assign n18488 = n18486 | n18487 ;
  assign n18489 = n12724 | n18488 ;
  assign n31296 = ~n18489 ;
  assign n18490 = x[11] & n31296 ;
  assign n18491 = n27892 & n18489 ;
  assign n18492 = n18490 | n18491 ;
  assign n31297 = ~n18492 ;
  assign n18493 = n18485 & n31297 ;
  assign n31298 = ~n18485 ;
  assign n18495 = n31298 & n18492 ;
  assign n18496 = n18493 | n18495 ;
  assign n15344 = n5417 & n15308 ;
  assign n15284 = x[121] & n15246 ;
  assign n17319 = x[122] & n16288 ;
  assign n18497 = n15284 | n17319 ;
  assign n18498 = x[123] & n15244 ;
  assign n18499 = n18497 | n18498 ;
  assign n18500 = n15344 | n18499 ;
  assign n31299 = ~n18500 ;
  assign n18501 = x[8] & n31299 ;
  assign n18502 = n27845 & n18500 ;
  assign n18503 = n18501 | n18502 ;
  assign n31300 = ~n18503 ;
  assign n18504 = n18496 & n31300 ;
  assign n31301 = ~n18496 ;
  assign n18595 = n31301 & n18503 ;
  assign n18596 = n18504 | n18595 ;
  assign n19593 = n19589 & n19591 ;
  assign n19594 = n18606 | n19593 ;
  assign n31302 = ~n19594 ;
  assign n19595 = n18596 & n31302 ;
  assign n31303 = ~n18596 ;
  assign n19597 = n31303 & n19594 ;
  assign n19598 = n19595 | n19597 ;
  assign n18429 = n5388 & n18392 ;
  assign n18388 = x[124] & n18329 ;
  assign n18559 = x[125] & n18514 ;
  assign n19599 = n18388 | n18559 ;
  assign n19600 = x[126] & n18327 ;
  assign n19601 = n19599 | n19600 ;
  assign n19602 = n18429 | n19601 ;
  assign n19603 = x[5] | n19602 ;
  assign n19604 = x[5] & n19602 ;
  assign n31304 = ~n19604 ;
  assign n19605 = n19603 & n31304 ;
  assign n19606 = n19598 & n19605 ;
  assign n19793 = n19598 | n19605 ;
  assign n31305 = ~n19606 ;
  assign n19794 = n31305 & n19793 ;
  assign n19640 = n19631 & n19638 ;
  assign n19652 = n19640 | n19651 ;
  assign n19684 = n5360 & n19656 ;
  assign n19728 = x[127] & n19723 ;
  assign n19788 = n19684 | n19728 ;
  assign n31306 = ~n19788 ;
  assign n19789 = x[2] & n31306 ;
  assign n19790 = n27790 & n19684 ;
  assign n19791 = n19789 | n19790 ;
  assign n19792 = n19652 & n19791 ;
  assign n19795 = n19652 | n19791 ;
  assign n31307 = ~n19792 ;
  assign n19796 = n31307 & n19795 ;
  assign n19797 = n19794 & n19796 ;
  assign n19802 = n19794 | n19796 ;
  assign n31308 = ~n19797 ;
  assign n19803 = n31308 & n19802 ;
  assign n19828 = n19825 & n19826 ;
  assign n19901 = n19828 | n19900 ;
  assign n31309 = ~n19901 ;
  assign n19902 = n19803 & n31309 ;
  assign n31310 = ~n19803 ;
  assign n19904 = n31310 & n19901 ;
  assign n19905 = n19902 | n19904 ;
  assign n23113 = n19948 | n23112 ;
  assign n23114 = n19905 | n23113 ;
  assign n23115 = n19905 & n23113 ;
  assign n31311 = ~n23115 ;
  assign n194 = n23114 & n31311 ;
  assign n19596 = n18596 & n19594 ;
  assign n19607 = n19596 | n19606 ;
  assign n18424 = n5629 & n18392 ;
  assign n18342 = x[125] & n18329 ;
  assign n18546 = x[126] & n18514 ;
  assign n19608 = n18342 | n18546 ;
  assign n19609 = x[127] & n18327 ;
  assign n19610 = n19608 | n19609 ;
  assign n19611 = n18424 | n19610 ;
  assign n31312 = ~n19611 ;
  assign n19612 = x[5] & n31312 ;
  assign n19613 = n27813 & n19611 ;
  assign n19614 = n19612 | n19613 ;
  assign n19615 = n19607 | n19614 ;
  assign n19616 = n19607 & n19614 ;
  assign n31313 = ~n19616 ;
  assign n19617 = n19615 & n31313 ;
  assign n12730 = n4985 & n12695 ;
  assign n12690 = x[119] & n12633 ;
  assign n14379 = x[120] & n13533 ;
  assign n17352 = n12690 | n14379 ;
  assign n17353 = x[121] & n12631 ;
  assign n17354 = n17352 | n17353 ;
  assign n17355 = n12730 | n17354 ;
  assign n31314 = ~n17355 ;
  assign n17356 = x[11] & n31314 ;
  assign n17357 = n27892 & n17355 ;
  assign n17358 = n17356 | n17357 ;
  assign n18296 = n17368 | n18295 ;
  assign n18297 = n17358 | n18296 ;
  assign n18298 = n17358 & n18296 ;
  assign n31315 = ~n18298 ;
  assign n18299 = n18297 & n31315 ;
  assign n8741 = n4474 & n8706 ;
  assign n8666 = x[113] & n8645 ;
  assign n9874 = x[114] & n9278 ;
  assign n15411 = n8666 | n9874 ;
  assign n15412 = x[115] & n8643 ;
  assign n15413 = n15411 | n15412 ;
  assign n15414 = n8741 | n15413 ;
  assign n31316 = ~n15414 ;
  assign n15415 = x[17] & n31316 ;
  assign n15416 = n28039 & n15414 ;
  assign n15417 = n15415 | n15416 ;
  assign n15428 = n15424 & n15426 ;
  assign n16254 = n16250 & n16252 ;
  assign n16255 = n15428 | n16254 ;
  assign n16256 = n15417 | n16255 ;
  assign n16257 = n15417 & n16255 ;
  assign n31317 = ~n16257 ;
  assign n16258 = n16256 & n31317 ;
  assign n7212 = n4442 & n7162 ;
  assign n7150 = x[110] & n7100 ;
  assign n7727 = x[111] & n7647 ;
  assign n14460 = n7150 | n7727 ;
  assign n14461 = x[112] & n7098 ;
  assign n14462 = n14460 | n14461 ;
  assign n14463 = n7212 | n14462 ;
  assign n31318 = ~n14463 ;
  assign n14464 = x[20] & n31318 ;
  assign n14465 = n28114 & n14463 ;
  assign n14466 = n14464 | n14465 ;
  assign n14479 = n14470 & n14477 ;
  assign n15196 = n14481 & n15194 ;
  assign n15197 = n14479 | n15196 ;
  assign n15198 = n14466 | n15197 ;
  assign n15199 = n14466 & n15197 ;
  assign n31319 = ~n15199 ;
  assign n15200 = n15198 & n31319 ;
  assign n5349 = n3639 & n5302 ;
  assign n5291 = x[107] & n5240 ;
  assign n6272 = x[108] & n6179 ;
  assign n14257 = n5291 | n6272 ;
  assign n14258 = x[109] & n5238 ;
  assign n14259 = n14257 | n14258 ;
  assign n14260 = n5349 | n14259 ;
  assign n31320 = ~n14260 ;
  assign n14261 = x[23] & n31320 ;
  assign n14262 = n28221 & n14260 ;
  assign n14263 = n14261 | n14262 ;
  assign n31321 = ~n14263 ;
  assign n14264 = n14256 & n31321 ;
  assign n14265 = n31281 & n14263 ;
  assign n14266 = n14264 | n14265 ;
  assign n3227 = n452 & n3223 ;
  assign n361 = x[104] & n330 ;
  assign n423 = x[105] & n390 ;
  assign n12812 = n361 | n423 ;
  assign n12813 = x[106] & n322 ;
  assign n12814 = n12812 | n12813 ;
  assign n12815 = n3227 | n12814 ;
  assign n12816 = x[26] | n12815 ;
  assign n12817 = x[26] & n12815 ;
  assign n31322 = ~n12817 ;
  assign n12818 = n12816 & n31322 ;
  assign n12828 = n12819 & n12826 ;
  assign n13466 = n12830 & n13464 ;
  assign n13467 = n12828 | n13466 ;
  assign n31323 = ~n13467 ;
  assign n13468 = n12818 & n31323 ;
  assign n31324 = ~n12818 ;
  assign n13470 = n31324 & n13467 ;
  assign n13471 = n13468 | n13470 ;
  assign n12548 = n12012 | n12547 ;
  assign n4510 = x[103] & n4504 ;
  assign n12549 = x[101] & n4514 ;
  assign n12550 = x[102] & n4572 ;
  assign n12551 = n12549 | n12550 ;
  assign n12552 = n4510 | n12551 ;
  assign n12553 = n2626 & n4632 ;
  assign n12554 = n12552 | n12553 ;
  assign n12555 = n28483 & n12554 ;
  assign n31325 = ~n12554 ;
  assign n12556 = x[29] & n31325 ;
  assign n12557 = n12555 | n12556 ;
  assign n31326 = ~n12557 ;
  assign n12558 = n12548 & n31326 ;
  assign n31327 = ~n12548 ;
  assign n12560 = n31327 & n12557 ;
  assign n12561 = n12558 | n12560 ;
  assign n4067 = n2438 & n4041 ;
  assign n3930 = x[95] & n3910 ;
  assign n4018 = x[96] & n3975 ;
  assign n11122 = n3930 | n4018 ;
  assign n11123 = x[97] & n3906 ;
  assign n11124 = n11122 | n11123 ;
  assign n11125 = n4067 | n11124 ;
  assign n31328 = ~n11125 ;
  assign n11126 = x[35] & n31328 ;
  assign n11127 = n28822 & n11125 ;
  assign n11128 = n11126 | n11127 ;
  assign n2657 = n1720 & n2635 ;
  assign n2543 = x[86] & n2492 ;
  assign n2594 = x[87] & n2557 ;
  assign n9129 = n2543 | n2594 ;
  assign n9130 = x[88] & n2488 ;
  assign n9131 = n9129 | n9130 ;
  assign n9132 = n2657 | n9131 ;
  assign n9133 = x[44] | n9132 ;
  assign n9134 = x[44] & n9132 ;
  assign n31329 = ~n9134 ;
  assign n9135 = n9133 & n31329 ;
  assign n1746 = n1690 & n1741 ;
  assign n1607 = x[77] & n1551 ;
  assign n1650 = x[78] & n1616 ;
  assign n7470 = n1607 | n1650 ;
  assign n7471 = x[79] & n1547 ;
  assign n7472 = n7470 | n7471 ;
  assign n7473 = n1746 | n7472 ;
  assign n7474 = x[53] | n7473 ;
  assign n7475 = x[53] & n7473 ;
  assign n31330 = ~n7475 ;
  assign n7476 = n7474 & n31330 ;
  assign n7465 = n7461 & n7463 ;
  assign n7466 = n7462 | n7465 ;
  assign n6521 = n6399 | n6520 ;
  assign n27783 = x[66] & n27215 ;
  assign n836 = x[67] & n805 ;
  assign n5965 = n27783 | n836 ;
  assign n5966 = x[2] | n5965 ;
  assign n5967 = x[2] & n5965 ;
  assign n31331 = ~n5967 ;
  assign n5968 = n5966 & n31331 ;
  assign n885 = x[70] & n881 ;
  assign n5969 = x[68] & n900 ;
  assign n5970 = x[69] & n949 ;
  assign n5971 = n5969 | n5970 ;
  assign n5972 = n885 | n5971 ;
  assign n5990 = n1006 & n5976 ;
  assign n5991 = n5972 | n5990 ;
  assign n5992 = n30886 & n5991 ;
  assign n31332 = ~n5991 ;
  assign n5993 = x[62] & n31332 ;
  assign n5994 = n5992 | n5993 ;
  assign n31333 = ~n5994 ;
  assign n5995 = n5968 & n31333 ;
  assign n31334 = ~n5968 ;
  assign n6522 = n31334 & n5994 ;
  assign n6523 = n5995 | n6522 ;
  assign n6524 = n6521 & n6523 ;
  assign n6525 = n6521 | n6523 ;
  assign n31335 = ~n6524 ;
  assign n6526 = n31335 & n6525 ;
  assign n3742 = n1217 & n3733 ;
  assign n1133 = x[71] & n1079 ;
  assign n1199 = x[72] & n1144 ;
  assign n6527 = n1133 | n1199 ;
  assign n6528 = x[73] & n1075 ;
  assign n6529 = n6527 | n6528 ;
  assign n6530 = n3742 | n6529 ;
  assign n31336 = ~n6530 ;
  assign n6531 = x[59] & n31336 ;
  assign n6532 = n30638 & n6530 ;
  assign n6533 = n6531 | n6532 ;
  assign n31337 = ~n6533 ;
  assign n6534 = n6526 & n31337 ;
  assign n31338 = ~n6526 ;
  assign n6904 = n31338 & n6533 ;
  assign n6905 = n6534 | n6904 ;
  assign n31339 = ~n6905 ;
  assign n6906 = n6903 & n31339 ;
  assign n6907 = n31237 & n6905 ;
  assign n6908 = n6906 | n6907 ;
  assign n2757 = n1457 & n2750 ;
  assign n1379 = x[74] & n1319 ;
  assign n1420 = x[75] & n1384 ;
  assign n6909 = n1379 | n1420 ;
  assign n6910 = x[76] & n1315 ;
  assign n6911 = n6909 | n6910 ;
  assign n6912 = n2757 | n6911 ;
  assign n31340 = ~n6912 ;
  assign n6913 = x[56] & n31340 ;
  assign n6914 = n30379 & n6912 ;
  assign n6915 = n6913 | n6914 ;
  assign n31341 = ~n6915 ;
  assign n6916 = n6908 & n31341 ;
  assign n31342 = ~n6908 ;
  assign n7467 = n31342 & n6915 ;
  assign n7468 = n6916 | n7467 ;
  assign n7469 = n7466 & n7468 ;
  assign n7477 = n7466 | n7468 ;
  assign n31343 = ~n7469 ;
  assign n7478 = n31343 & n7477 ;
  assign n7479 = n7476 & n7478 ;
  assign n7790 = n7476 | n7478 ;
  assign n31344 = ~n7479 ;
  assign n7791 = n31344 & n7790 ;
  assign n7991 = n7987 & n7989 ;
  assign n7992 = n7801 | n7991 ;
  assign n31345 = ~n7992 ;
  assign n7993 = n7791 & n31345 ;
  assign n31346 = ~n7791 ;
  assign n7995 = n31346 & n7992 ;
  assign n7996 = n7993 | n7995 ;
  assign n2019 = n1003 & n2007 ;
  assign n1901 = x[80] & n1866 ;
  assign n1988 = x[81] & n1931 ;
  assign n7997 = n1901 | n1988 ;
  assign n7998 = x[82] & n1862 ;
  assign n7999 = n7997 | n7998 ;
  assign n8000 = n2019 | n7999 ;
  assign n31347 = ~n8000 ;
  assign n8001 = x[50] & n31347 ;
  assign n8002 = n29865 & n8000 ;
  assign n8003 = n8001 | n8002 ;
  assign n31348 = ~n8003 ;
  assign n8004 = n7996 & n31348 ;
  assign n31349 = ~n7996 ;
  assign n8242 = n31349 & n8003 ;
  assign n8243 = n8004 | n8242 ;
  assign n8486 = n8254 | n8485 ;
  assign n31350 = ~n8486 ;
  assign n8487 = n8243 & n31350 ;
  assign n31351 = ~n8243 ;
  assign n8489 = n31351 & n8486 ;
  assign n8490 = n8487 | n8489 ;
  assign n2340 = n1239 & n2321 ;
  assign n2208 = x[83] & n2179 ;
  assign n2298 = x[84] & n2244 ;
  assign n8491 = n2208 | n2298 ;
  assign n8492 = x[85] & n2175 ;
  assign n8493 = n8491 | n8492 ;
  assign n8494 = n2340 | n8493 ;
  assign n31352 = ~n8494 ;
  assign n8495 = x[47] & n31352 ;
  assign n8496 = n29621 & n8494 ;
  assign n8497 = n8495 | n8496 ;
  assign n31353 = ~n8497 ;
  assign n8498 = n8490 & n31353 ;
  assign n31354 = ~n8490 ;
  assign n8836 = n31354 & n8497 ;
  assign n8837 = n8498 | n8836 ;
  assign n8848 = n8839 & n8846 ;
  assign n9124 = n9121 & n9123 ;
  assign n9126 = n8848 | n9124 ;
  assign n31355 = ~n9126 ;
  assign n9127 = n8837 & n31355 ;
  assign n31356 = ~n8837 ;
  assign n9136 = n31356 & n9126 ;
  assign n9137 = n9127 | n9136 ;
  assign n9138 = n9135 & n9137 ;
  assign n9329 = n9135 | n9137 ;
  assign n31357 = ~n9138 ;
  assign n9330 = n31357 & n9329 ;
  assign n9672 = n9341 | n9671 ;
  assign n31358 = ~n9672 ;
  assign n9673 = n9330 & n31358 ;
  assign n31359 = ~n9330 ;
  assign n9675 = n31359 & n9672 ;
  assign n9676 = n9673 | n9675 ;
  assign n3166 = n2046 & n3162 ;
  assign n3083 = x[89] & n3031 ;
  assign n3152 = x[90] & n3096 ;
  assign n9677 = n3083 | n3152 ;
  assign n9678 = x[91] & n3027 ;
  assign n9679 = n9677 | n9678 ;
  assign n9680 = n3166 | n9679 ;
  assign n31360 = ~n9680 ;
  assign n9681 = x[41] & n31360 ;
  assign n9682 = n29184 & n9680 ;
  assign n9683 = n9681 | n9682 ;
  assign n31361 = ~n9683 ;
  assign n9684 = n9676 & n31361 ;
  assign n31362 = ~n9676 ;
  assign n9980 = n31362 & n9683 ;
  assign n9981 = n9684 | n9980 ;
  assign n9992 = n9983 & n9990 ;
  assign n10362 = n9994 & n10360 ;
  assign n10363 = n9992 | n10362 ;
  assign n10364 = n9981 | n10363 ;
  assign n10365 = n9981 & n10363 ;
  assign n31363 = ~n10365 ;
  assign n10366 = n10364 & n31363 ;
  assign n3609 = n2410 & n3574 ;
  assign n3488 = x[92] & n3443 ;
  assign n3511 = x[93] & n3508 ;
  assign n10367 = n3488 | n3511 ;
  assign n10368 = x[94] & n3439 ;
  assign n10369 = n10367 | n10368 ;
  assign n10370 = n3609 | n10369 ;
  assign n31364 = ~n10370 ;
  assign n10371 = x[38] & n31364 ;
  assign n10372 = n28996 & n10370 ;
  assign n10373 = n10371 | n10372 ;
  assign n31365 = ~n10373 ;
  assign n10374 = n10366 & n31365 ;
  assign n31366 = ~n10366 ;
  assign n10662 = n31366 & n10373 ;
  assign n10663 = n10374 | n10662 ;
  assign n10674 = n10665 & n10672 ;
  assign n11119 = n10676 & n11117 ;
  assign n11120 = n10674 | n11119 ;
  assign n11121 = n10663 | n11120 ;
  assign n11129 = n10663 & n11120 ;
  assign n31367 = ~n11129 ;
  assign n11130 = n11121 & n31367 ;
  assign n11131 = n11128 & n11130 ;
  assign n11733 = n11128 | n11130 ;
  assign n31368 = ~n11131 ;
  assign n11734 = n31368 & n11733 ;
  assign n658 = x[100] & n652 ;
  assign n11723 = x[98] & n663 ;
  assign n11724 = x[99] & n720 ;
  assign n11725 = n11723 | n11724 ;
  assign n11726 = n658 | n11725 ;
  assign n11727 = n779 & n2466 ;
  assign n11728 = n11726 | n11727 ;
  assign n11729 = n28658 & n11728 ;
  assign n31369 = ~n11728 ;
  assign n11730 = x[32] & n31369 ;
  assign n11731 = n11729 | n11730 ;
  assign n11732 = n11721 | n11731 ;
  assign n11735 = n11721 & n11731 ;
  assign n31370 = ~n11735 ;
  assign n11736 = n11732 & n31370 ;
  assign n31371 = ~n11736 ;
  assign n11737 = n11734 & n31371 ;
  assign n31372 = ~n11734 ;
  assign n12562 = n31372 & n11736 ;
  assign n12563 = n11737 | n12562 ;
  assign n31373 = ~n12563 ;
  assign n12564 = n12561 & n31373 ;
  assign n31374 = ~n12561 ;
  assign n13472 = n31374 & n12563 ;
  assign n13473 = n12564 | n13472 ;
  assign n13474 = n13471 & n13473 ;
  assign n14267 = n13471 | n13473 ;
  assign n14268 = n14266 & n14267 ;
  assign n31375 = ~n13474 ;
  assign n14269 = n31375 & n14268 ;
  assign n31376 = ~n14269 ;
  assign n14270 = n14266 & n31376 ;
  assign n15201 = n14267 & n31376 ;
  assign n15202 = n31375 & n15201 ;
  assign n15203 = n14270 | n15202 ;
  assign n15204 = n15200 & n15203 ;
  assign n16260 = n15200 | n15203 ;
  assign n16261 = n16258 & n16260 ;
  assign n31377 = ~n15204 ;
  assign n16262 = n31377 & n16261 ;
  assign n31378 = ~n16262 ;
  assign n16263 = n16258 & n31378 ;
  assign n16259 = n31377 & n16258 ;
  assign n31379 = ~n16259 ;
  assign n17230 = n31379 & n16260 ;
  assign n17231 = n31377 & n17230 ;
  assign n17232 = n16263 | n17231 ;
  assign n17218 = n17215 | n17217 ;
  assign n11852 = x[118] & n10479 ;
  assign n17219 = x[116] & n10481 ;
  assign n17220 = x[117] & n11232 ;
  assign n17221 = n17219 | n17220 ;
  assign n17222 = n11852 | n17221 ;
  assign n17223 = n784 & n10542 ;
  assign n17224 = n17222 | n17223 ;
  assign n17225 = n27956 & n17224 ;
  assign n31380 = ~n17224 ;
  assign n17226 = x[14] & n31380 ;
  assign n17227 = n17225 | n17226 ;
  assign n31381 = ~n17227 ;
  assign n17228 = n17218 & n31381 ;
  assign n31382 = ~n17218 ;
  assign n17233 = n31382 & n17227 ;
  assign n17234 = n17228 | n17233 ;
  assign n17235 = n17232 | n17234 ;
  assign n17236 = n17232 & n17234 ;
  assign n31383 = ~n17236 ;
  assign n18300 = n17235 & n31383 ;
  assign n18301 = n18299 | n18300 ;
  assign n18302 = n18299 & n18300 ;
  assign n31384 = ~n18302 ;
  assign n18509 = n18301 & n31384 ;
  assign n15311 = n5838 & n15308 ;
  assign n15267 = x[122] & n15246 ;
  assign n17311 = x[123] & n16288 ;
  assign n18477 = n15267 | n17311 ;
  assign n18478 = x[124] & n15244 ;
  assign n18479 = n18477 | n18478 ;
  assign n18480 = n15311 | n18479 ;
  assign n18481 = x[8] | n18480 ;
  assign n18482 = x[8] & n18480 ;
  assign n31385 = ~n18482 ;
  assign n18483 = n18481 & n31385 ;
  assign n18494 = n18485 & n18492 ;
  assign n18505 = n18496 & n18503 ;
  assign n18506 = n18494 | n18505 ;
  assign n31386 = ~n18506 ;
  assign n18507 = n18483 & n31386 ;
  assign n31387 = ~n18483 ;
  assign n18510 = n31387 & n18506 ;
  assign n18511 = n18507 | n18510 ;
  assign n18512 = n18509 & n18511 ;
  assign n19618 = n18509 | n18511 ;
  assign n31388 = ~n18512 ;
  assign n19619 = n31388 & n19618 ;
  assign n19620 = n19617 | n19619 ;
  assign n19621 = n19617 & n19619 ;
  assign n31389 = ~n19621 ;
  assign n19629 = n19620 & n31389 ;
  assign n19798 = n19792 | n19797 ;
  assign n19799 = n19629 | n19798 ;
  assign n19800 = n19629 & n19798 ;
  assign n31390 = ~n19800 ;
  assign n19801 = n19799 & n31390 ;
  assign n19903 = n19803 & n19901 ;
  assign n23116 = n19903 | n23115 ;
  assign n23117 = n19801 & n23116 ;
  assign n27724 = n19801 | n23116 ;
  assign n31391 = ~n23117 ;
  assign n195 = n31391 & n27724 ;
  assign n23118 = n19800 | n23117 ;
  assign n19622 = n19616 | n19621 ;
  assign n10581 = n5047 & n10542 ;
  assign n10530 = x[117] & n10481 ;
  assign n11898 = x[118] & n11232 ;
  assign n15404 = n10530 | n11898 ;
  assign n15405 = x[119] & n10479 ;
  assign n15406 = n15404 | n15405 ;
  assign n15407 = n10581 | n15406 ;
  assign n31392 = ~n15407 ;
  assign n15408 = x[14] & n31392 ;
  assign n15409 = n27956 & n15407 ;
  assign n15410 = n15408 | n15409 ;
  assign n16264 = n16257 | n16262 ;
  assign n16265 = n15410 | n16264 ;
  assign n16266 = n15410 & n16264 ;
  assign n31393 = ~n16266 ;
  assign n16267 = n16265 & n31393 ;
  assign n7211 = n4087 & n7162 ;
  assign n7148 = x[111] & n7100 ;
  assign n7704 = x[112] & n7647 ;
  assign n13553 = n7148 | n7704 ;
  assign n13554 = x[113] & n7098 ;
  assign n13555 = n13553 | n13554 ;
  assign n13556 = n7211 | n13555 ;
  assign n31394 = ~n13556 ;
  assign n13557 = x[20] & n31394 ;
  assign n13558 = n28114 & n13556 ;
  assign n13559 = n13557 | n13558 ;
  assign n14271 = n14256 & n14263 ;
  assign n14272 = n14269 | n14271 ;
  assign n14273 = n13559 | n14272 ;
  assign n14274 = n13559 & n14272 ;
  assign n31395 = ~n14274 ;
  assign n14275 = n14273 & n31395 ;
  assign n3204 = n452 & n3199 ;
  assign n381 = x[105] & n330 ;
  assign n400 = x[106] & n390 ;
  assign n11994 = n381 | n400 ;
  assign n11995 = x[107] & n322 ;
  assign n11996 = n11994 | n11995 ;
  assign n11997 = n3204 | n11996 ;
  assign n11998 = x[26] | n11997 ;
  assign n11999 = x[26] & n11997 ;
  assign n31396 = ~n11999 ;
  assign n12000 = n11998 & n31396 ;
  assign n12559 = n12548 & n12557 ;
  assign n12565 = n12561 & n12563 ;
  assign n12566 = n12559 | n12565 ;
  assign n31397 = ~n12566 ;
  assign n12567 = n12000 & n31397 ;
  assign n31398 = ~n12000 ;
  assign n12569 = n31398 & n12566 ;
  assign n12570 = n12567 | n12569 ;
  assign n11132 = n11129 | n11131 ;
  assign n655 = x[101] & n652 ;
  assign n11133 = x[99] & n663 ;
  assign n11134 = x[100] & n720 ;
  assign n11135 = n11133 | n11134 ;
  assign n11136 = n655 | n11135 ;
  assign n11137 = n779 & n2977 ;
  assign n11138 = n11136 | n11137 ;
  assign n11139 = n28658 & n11138 ;
  assign n31399 = ~n11138 ;
  assign n11140 = x[32] & n31399 ;
  assign n11141 = n11139 | n11140 ;
  assign n31400 = ~n11141 ;
  assign n11142 = n11132 & n31400 ;
  assign n31401 = ~n11132 ;
  assign n11144 = n31401 & n11141 ;
  assign n11145 = n11142 | n11144 ;
  assign n4073 = n2841 & n4041 ;
  assign n3942 = x[96] & n3910 ;
  assign n4034 = x[97] & n3975 ;
  assign n10381 = n3942 | n4034 ;
  assign n10382 = x[98] & n3906 ;
  assign n10383 = n10381 | n10382 ;
  assign n10384 = n4073 | n10383 ;
  assign n10385 = x[35] | n10384 ;
  assign n10386 = x[35] & n10384 ;
  assign n31402 = ~n10386 ;
  assign n10387 = n10385 & n31402 ;
  assign n10375 = n10366 & n10373 ;
  assign n10376 = n10365 | n10375 ;
  assign n1702 = n1270 & n1690 ;
  assign n1568 = x[78] & n1551 ;
  assign n1672 = x[79] & n1616 ;
  assign n6922 = n1568 | n1672 ;
  assign n6923 = x[80] & n1547 ;
  assign n6924 = n6922 | n6923 ;
  assign n6925 = n1702 | n6924 ;
  assign n6926 = x[53] | n6925 ;
  assign n6927 = x[53] & n6925 ;
  assign n31403 = ~n6927 ;
  assign n6928 = n6926 & n31403 ;
  assign n925 = x[69] & n900 ;
  assign n967 = x[70] & n949 ;
  assign n4787 = n925 | n967 ;
  assign n4788 = x[71] & n881 ;
  assign n4789 = n4787 | n4788 ;
  assign n4802 = n1006 & n4790 ;
  assign n4804 = n4789 | n4802 ;
  assign n4805 = x[62] | n4804 ;
  assign n4806 = x[62] & n4804 ;
  assign n31404 = ~n4806 ;
  assign n4807 = n4805 & n31404 ;
  assign n27764 = x[67] & n27215 ;
  assign n851 = x[68] & n805 ;
  assign n4784 = n27764 | n851 ;
  assign n31405 = ~n4784 ;
  assign n4785 = x[2] & n31405 ;
  assign n4808 = n27790 & n4784 ;
  assign n4809 = n4785 | n4808 ;
  assign n31406 = ~n4809 ;
  assign n4810 = n4807 & n31406 ;
  assign n31407 = ~n4807 ;
  assign n5963 = n31407 & n4809 ;
  assign n5964 = n4810 | n5963 ;
  assign n5996 = n5968 & n5994 ;
  assign n5997 = n5967 | n5996 ;
  assign n31408 = ~n5997 ;
  assign n5998 = n5964 & n31408 ;
  assign n31409 = ~n5964 ;
  assign n6000 = n31409 & n5997 ;
  assign n6001 = n5998 | n6000 ;
  assign n2726 = n1217 & n2722 ;
  assign n1140 = x[72] & n1079 ;
  assign n1155 = x[73] & n1144 ;
  assign n6002 = n1140 | n1155 ;
  assign n6003 = x[74] & n1075 ;
  assign n6004 = n6002 | n6003 ;
  assign n6005 = n2726 | n6004 ;
  assign n31410 = ~n6005 ;
  assign n6006 = x[59] & n31410 ;
  assign n6007 = n30638 & n6005 ;
  assign n6008 = n6006 | n6007 ;
  assign n31411 = ~n6008 ;
  assign n6009 = n6001 & n31411 ;
  assign n31412 = ~n6001 ;
  assign n6373 = n31412 & n6008 ;
  assign n6374 = n6009 | n6373 ;
  assign n6535 = n6526 & n6533 ;
  assign n6536 = n6524 | n6535 ;
  assign n31413 = ~n6536 ;
  assign n6537 = n6374 & n31413 ;
  assign n31414 = ~n6374 ;
  assign n6539 = n31414 & n6536 ;
  assign n6540 = n6537 | n6539 ;
  assign n1779 = n1457 & n1775 ;
  assign n1362 = x[75] & n1319 ;
  assign n1435 = x[76] & n1384 ;
  assign n6541 = n1362 | n1435 ;
  assign n6542 = x[77] & n1315 ;
  assign n6543 = n6541 | n6542 ;
  assign n6544 = n1779 | n6543 ;
  assign n31415 = ~n6544 ;
  assign n6545 = x[56] & n31415 ;
  assign n6546 = n30379 & n6544 ;
  assign n6547 = n6545 | n6546 ;
  assign n31416 = ~n6547 ;
  assign n6548 = n6540 & n31416 ;
  assign n31417 = ~n6540 ;
  assign n6796 = n31417 & n6547 ;
  assign n6797 = n6548 | n6796 ;
  assign n6917 = n6908 & n6915 ;
  assign n6918 = n6903 & n6905 ;
  assign n6919 = n6917 | n6918 ;
  assign n6920 = n6797 | n6919 ;
  assign n6921 = n6797 & n6919 ;
  assign n31418 = ~n6921 ;
  assign n6929 = n6920 & n31418 ;
  assign n6930 = n6928 & n6929 ;
  assign n7307 = n6928 | n6929 ;
  assign n31419 = ~n6930 ;
  assign n7308 = n31419 & n7307 ;
  assign n7480 = n7469 | n7479 ;
  assign n31420 = ~n7480 ;
  assign n7481 = n7308 & n31420 ;
  assign n31421 = ~n7308 ;
  assign n7483 = n31421 & n7480 ;
  assign n7484 = n7481 | n7483 ;
  assign n2015 = n1057 & n2007 ;
  assign n1925 = x[81] & n1866 ;
  assign n1945 = x[82] & n1931 ;
  assign n7485 = n1925 | n1945 ;
  assign n7486 = x[83] & n1862 ;
  assign n7487 = n7485 | n7486 ;
  assign n7488 = n2015 | n7487 ;
  assign n31422 = ~n7488 ;
  assign n7489 = x[50] & n31422 ;
  assign n7490 = n29865 & n7488 ;
  assign n7491 = n7489 | n7490 ;
  assign n31423 = ~n7491 ;
  assign n7492 = n7484 & n31423 ;
  assign n31424 = ~n7484 ;
  assign n7788 = n31424 & n7491 ;
  assign n7789 = n7492 | n7788 ;
  assign n7994 = n7791 & n7992 ;
  assign n8005 = n7996 & n8003 ;
  assign n8006 = n7994 | n8005 ;
  assign n31425 = ~n8006 ;
  assign n8007 = n7789 & n31425 ;
  assign n31426 = ~n7789 ;
  assign n8009 = n31426 & n8006 ;
  assign n8010 = n8007 | n8009 ;
  assign n2325 = n1213 & n2321 ;
  assign n2222 = x[84] & n2179 ;
  assign n2296 = x[85] & n2244 ;
  assign n8011 = n2222 | n2296 ;
  assign n8012 = x[86] & n2175 ;
  assign n8013 = n8011 | n8012 ;
  assign n8014 = n2325 | n8013 ;
  assign n31427 = ~n8014 ;
  assign n8015 = x[47] & n31427 ;
  assign n8016 = n29621 & n8014 ;
  assign n8017 = n8015 | n8016 ;
  assign n31428 = ~n8017 ;
  assign n8018 = n8010 & n31428 ;
  assign n31429 = ~n8010 ;
  assign n8240 = n31429 & n8017 ;
  assign n8241 = n8018 | n8240 ;
  assign n8488 = n8243 & n8486 ;
  assign n8499 = n8490 & n8497 ;
  assign n8500 = n8488 | n8499 ;
  assign n31430 = ~n8500 ;
  assign n8501 = n8241 & n31430 ;
  assign n31431 = ~n8241 ;
  assign n8503 = n31431 & n8500 ;
  assign n8504 = n8501 | n8503 ;
  assign n2654 = n1453 & n2635 ;
  assign n2549 = x[87] & n2492 ;
  assign n2602 = x[88] & n2557 ;
  assign n8505 = n2549 | n2602 ;
  assign n8506 = x[89] & n2488 ;
  assign n8507 = n8505 | n8506 ;
  assign n8508 = n2654 | n8507 ;
  assign n31432 = ~n8508 ;
  assign n8509 = x[44] & n31432 ;
  assign n8510 = n29400 & n8508 ;
  assign n8511 = n8509 | n8510 ;
  assign n31433 = ~n8511 ;
  assign n8512 = n8504 & n31433 ;
  assign n31434 = ~n8504 ;
  assign n8834 = n31434 & n8511 ;
  assign n8835 = n8512 | n8834 ;
  assign n9128 = n8837 & n9126 ;
  assign n9139 = n9128 | n9138 ;
  assign n31435 = ~n9139 ;
  assign n9140 = n8835 & n31435 ;
  assign n31436 = ~n8835 ;
  assign n9142 = n31436 & n9139 ;
  assign n9143 = n9140 | n9142 ;
  assign n3183 = n1841 & n3162 ;
  assign n3089 = x[90] & n3031 ;
  assign n3153 = x[91] & n3096 ;
  assign n9144 = n3089 | n3153 ;
  assign n9145 = x[92] & n3027 ;
  assign n9146 = n9144 | n9145 ;
  assign n9147 = n3183 | n9146 ;
  assign n31437 = ~n9147 ;
  assign n9148 = x[41] & n31437 ;
  assign n9149 = n29184 & n9147 ;
  assign n9150 = n9148 | n9149 ;
  assign n31438 = ~n9150 ;
  assign n9151 = n9143 & n31438 ;
  assign n31439 = ~n9143 ;
  assign n9327 = n31439 & n9150 ;
  assign n9328 = n9151 | n9327 ;
  assign n9674 = n9330 & n9672 ;
  assign n9685 = n9676 & n9683 ;
  assign n9686 = n9674 | n9685 ;
  assign n31440 = ~n9686 ;
  assign n9687 = n9328 & n31440 ;
  assign n31441 = ~n9328 ;
  assign n9689 = n31441 & n9686 ;
  assign n9690 = n9687 | n9689 ;
  assign n3599 = n2152 & n3574 ;
  assign n3500 = x[93] & n3443 ;
  assign n3567 = x[94] & n3508 ;
  assign n9691 = n3500 | n3567 ;
  assign n9692 = x[95] & n3439 ;
  assign n9693 = n9691 | n9692 ;
  assign n9694 = n3599 | n9693 ;
  assign n31442 = ~n9694 ;
  assign n9695 = x[38] & n31442 ;
  assign n9696 = n28996 & n9694 ;
  assign n9697 = n9695 | n9696 ;
  assign n31443 = ~n9697 ;
  assign n9698 = n9690 & n31443 ;
  assign n31444 = ~n9690 ;
  assign n10377 = n31444 & n9697 ;
  assign n10378 = n9698 | n10377 ;
  assign n31445 = ~n10376 ;
  assign n10379 = n31445 & n10378 ;
  assign n31446 = ~n10378 ;
  assign n10388 = n10376 & n31446 ;
  assign n10389 = n10379 | n10388 ;
  assign n31447 = ~n10389 ;
  assign n10390 = n10387 & n31447 ;
  assign n31448 = ~n10387 ;
  assign n11146 = n31448 & n10389 ;
  assign n11147 = n10390 | n11146 ;
  assign n31449 = ~n11147 ;
  assign n11148 = n11145 & n31449 ;
  assign n31450 = ~n11145 ;
  assign n11751 = n31450 & n11147 ;
  assign n11752 = n11148 | n11751 ;
  assign n11738 = n11734 & n11736 ;
  assign n11739 = n11735 | n11738 ;
  assign n4508 = x[104] & n4504 ;
  assign n11740 = x[102] & n4514 ;
  assign n11741 = x[103] & n4572 ;
  assign n11742 = n11740 | n11741 ;
  assign n11743 = n4508 | n11742 ;
  assign n11744 = n3001 & n4632 ;
  assign n11745 = n11743 | n11744 ;
  assign n11746 = n28483 & n11745 ;
  assign n31451 = ~n11745 ;
  assign n11747 = x[29] & n31451 ;
  assign n11748 = n11746 | n11747 ;
  assign n31452 = ~n11748 ;
  assign n11749 = n11739 & n31452 ;
  assign n31453 = ~n11739 ;
  assign n11753 = n31453 & n11748 ;
  assign n11754 = n11749 | n11753 ;
  assign n31454 = ~n11754 ;
  assign n11755 = n11752 & n31454 ;
  assign n31455 = ~n11752 ;
  assign n12571 = n31455 & n11754 ;
  assign n12572 = n11755 | n12571 ;
  assign n31456 = ~n12572 ;
  assign n12573 = n12570 & n31456 ;
  assign n31457 = ~n12570 ;
  assign n13478 = n31457 & n12572 ;
  assign n13479 = n12573 | n13478 ;
  assign n5341 = n3615 & n5302 ;
  assign n5285 = x[108] & n5240 ;
  assign n6263 = x[109] & n6179 ;
  assign n12805 = n5285 | n6263 ;
  assign n12806 = x[110] & n5238 ;
  assign n12807 = n12805 | n12806 ;
  assign n12808 = n5341 | n12807 ;
  assign n12809 = x[23] | n12808 ;
  assign n12810 = x[23] & n12808 ;
  assign n31458 = ~n12810 ;
  assign n12811 = n12809 & n31458 ;
  assign n13469 = n12818 & n13467 ;
  assign n13475 = n13469 | n13474 ;
  assign n31459 = ~n13475 ;
  assign n13476 = n12811 & n31459 ;
  assign n31460 = ~n12811 ;
  assign n13480 = n31460 & n13475 ;
  assign n13481 = n13476 | n13480 ;
  assign n31461 = ~n13481 ;
  assign n13482 = n13479 & n31461 ;
  assign n31462 = ~n13479 ;
  assign n14276 = n31462 & n13481 ;
  assign n14277 = n13482 | n14276 ;
  assign n14278 = n14275 | n14277 ;
  assign n14279 = n14275 & n14277 ;
  assign n31463 = ~n14279 ;
  assign n15208 = n14278 & n31463 ;
  assign n8744 = n4702 & n8706 ;
  assign n8650 = x[114] & n8645 ;
  assign n9852 = x[115] & n9278 ;
  assign n14453 = n8650 | n9852 ;
  assign n14454 = x[116] & n8643 ;
  assign n14455 = n14453 | n14454 ;
  assign n14456 = n8744 | n14455 ;
  assign n31464 = ~n14456 ;
  assign n14457 = x[17] & n31464 ;
  assign n14458 = n28039 & n14456 ;
  assign n14459 = n14457 | n14458 ;
  assign n15205 = n15199 | n15204 ;
  assign n15206 = n14459 | n15205 ;
  assign n15207 = n14459 & n15205 ;
  assign n31465 = ~n15207 ;
  assign n15209 = n15206 & n31465 ;
  assign n31466 = ~n15209 ;
  assign n15210 = n15208 & n31466 ;
  assign n31467 = ~n15208 ;
  assign n16268 = n31467 & n15209 ;
  assign n16269 = n15210 | n16268 ;
  assign n16270 = n16267 & n16269 ;
  assign n17249 = n16267 | n16269 ;
  assign n31468 = ~n16270 ;
  assign n17250 = n31468 & n17249 ;
  assign n17229 = n17218 & n17227 ;
  assign n17237 = n17229 | n17236 ;
  assign n14332 = x[122] & n12631 ;
  assign n17238 = x[120] & n12633 ;
  assign n17239 = x[121] & n13533 ;
  assign n17240 = n17238 | n17239 ;
  assign n17241 = n14332 | n17240 ;
  assign n17242 = n5022 & n12695 ;
  assign n17243 = n17241 | n17242 ;
  assign n17244 = n27892 & n17243 ;
  assign n31469 = ~n17243 ;
  assign n17245 = x[11] & n31469 ;
  assign n17246 = n17244 | n17245 ;
  assign n31470 = ~n17246 ;
  assign n17247 = n17237 & n31470 ;
  assign n31471 = ~n17237 ;
  assign n17251 = n31471 & n17246 ;
  assign n17252 = n17247 | n17251 ;
  assign n17253 = n17250 & n17252 ;
  assign n18315 = n17250 | n17252 ;
  assign n31472 = ~n17253 ;
  assign n18316 = n31472 & n18315 ;
  assign n18303 = n18298 | n18302 ;
  assign n17256 = x[125] & n15244 ;
  assign n18304 = x[123] & n15246 ;
  assign n18305 = x[124] & n16288 ;
  assign n18306 = n18304 | n18305 ;
  assign n18307 = n17256 | n18306 ;
  assign n18308 = n642 & n15308 ;
  assign n18309 = n18307 | n18308 ;
  assign n18310 = n27845 & n18309 ;
  assign n31473 = ~n18309 ;
  assign n18311 = x[8] & n31473 ;
  assign n18312 = n18310 | n18311 ;
  assign n31474 = ~n18312 ;
  assign n18313 = n18303 & n31474 ;
  assign n31475 = ~n18303 ;
  assign n18317 = n31475 & n18312 ;
  assign n18318 = n18313 | n18317 ;
  assign n18319 = n18316 & n18318 ;
  assign n18586 = n18316 | n18318 ;
  assign n31476 = ~n18319 ;
  assign n18587 = n31476 & n18586 ;
  assign n18508 = n18483 & n18506 ;
  assign n18513 = n18508 | n18512 ;
  assign n18397 = n6186 & n18392 ;
  assign n18576 = x[126] & n18329 ;
  assign n18577 = x[127] & n18514 ;
  assign n18578 = n18576 | n18577 ;
  assign n18579 = n18397 | n18578 ;
  assign n31477 = ~n18579 ;
  assign n18580 = x[5] & n31477 ;
  assign n18581 = n27813 & n18579 ;
  assign n18582 = n18580 | n18581 ;
  assign n18584 = n18513 | n18582 ;
  assign n18585 = n18513 & n18582 ;
  assign n31478 = ~n18585 ;
  assign n18588 = n18584 & n31478 ;
  assign n18589 = n18587 & n18588 ;
  assign n31479 = ~n18582 ;
  assign n19623 = n18513 & n31479 ;
  assign n31480 = ~n18513 ;
  assign n18583 = n31480 & n18582 ;
  assign n19624 = n18583 | n18587 ;
  assign n19625 = n19623 | n19624 ;
  assign n31481 = ~n18589 ;
  assign n19626 = n31481 & n19625 ;
  assign n31482 = ~n19622 ;
  assign n19627 = n31482 & n19626 ;
  assign n31483 = ~n19626 ;
  assign n23119 = n19622 & n31483 ;
  assign n23120 = n19627 | n23119 ;
  assign n23121 = n23118 & n23120 ;
  assign n27726 = n19627 | n23118 ;
  assign n27727 = n23119 | n27726 ;
  assign n31484 = ~n23121 ;
  assign n196 = n31484 & n27727 ;
  assign n19628 = n19622 & n19626 ;
  assign n23122 = n19628 | n23121 ;
  assign n18590 = n18585 | n18589 ;
  assign n18314 = n18303 & n18312 ;
  assign n18320 = n18314 | n18319 ;
  assign n18369 = x[127] & n18329 ;
  assign n18431 = n5360 & n18392 ;
  assign n18458 = n18369 | n18431 ;
  assign n31485 = ~n18458 ;
  assign n18459 = x[5] & n31485 ;
  assign n18460 = n27813 & n18458 ;
  assign n18461 = n18459 | n18460 ;
  assign n18462 = n18320 | n18461 ;
  assign n18463 = n18320 & n18461 ;
  assign n31486 = ~n18463 ;
  assign n18464 = n18462 & n31486 ;
  assign n12742 = n5417 & n12695 ;
  assign n12672 = x[121] & n12633 ;
  assign n14384 = x[122] & n13533 ;
  assign n15397 = n12672 | n14384 ;
  assign n15398 = x[123] & n12631 ;
  assign n15399 = n15397 | n15398 ;
  assign n15400 = n12742 | n15399 ;
  assign n15401 = x[11] | n15400 ;
  assign n15402 = x[11] & n15400 ;
  assign n31487 = ~n15402 ;
  assign n15403 = n15401 & n31487 ;
  assign n16271 = n16266 | n16270 ;
  assign n31488 = ~n16271 ;
  assign n16272 = n15403 & n31488 ;
  assign n31489 = ~n15403 ;
  assign n16274 = n31489 & n16271 ;
  assign n16275 = n16272 | n16274 ;
  assign n10582 = n4678 & n10542 ;
  assign n10536 = x[118] & n10481 ;
  assign n11882 = x[119] & n11232 ;
  assign n14446 = n10536 | n11882 ;
  assign n14447 = x[120] & n10479 ;
  assign n14448 = n14446 | n14447 ;
  assign n14449 = n10582 | n14448 ;
  assign n14450 = x[14] | n14449 ;
  assign n14451 = x[14] & n14449 ;
  assign n31490 = ~n14451 ;
  assign n14452 = n14450 & n31490 ;
  assign n15211 = n15208 & n15209 ;
  assign n15212 = n15207 | n15211 ;
  assign n31491 = ~n15212 ;
  assign n15213 = n14452 & n31491 ;
  assign n31492 = ~n14452 ;
  assign n15215 = n31492 & n15212 ;
  assign n15216 = n15213 | n15215 ;
  assign n14280 = n14274 | n14279 ;
  assign n9823 = x[117] & n8643 ;
  assign n14281 = x[115] & n8645 ;
  assign n14282 = x[116] & n9278 ;
  assign n14283 = n14281 | n14282 ;
  assign n14284 = n9823 | n14283 ;
  assign n14285 = n797 & n8706 ;
  assign n14286 = n14284 | n14285 ;
  assign n14287 = n28039 & n14286 ;
  assign n31493 = ~n14286 ;
  assign n14288 = x[17] & n31493 ;
  assign n14289 = n14287 | n14288 ;
  assign n14290 = n14280 | n14289 ;
  assign n14291 = n14280 & n14289 ;
  assign n31494 = ~n14291 ;
  assign n14292 = n14290 & n31494 ;
  assign n7179 = n4276 & n7162 ;
  assign n7130 = x[112] & n7100 ;
  assign n7697 = x[113] & n7647 ;
  assign n12798 = n7130 | n7697 ;
  assign n12799 = x[114] & n7098 ;
  assign n12800 = n12798 | n12799 ;
  assign n12801 = n7179 | n12800 ;
  assign n12802 = x[20] | n12801 ;
  assign n12803 = x[20] & n12801 ;
  assign n31495 = ~n12803 ;
  assign n12804 = n12802 & n31495 ;
  assign n13477 = n12811 & n13475 ;
  assign n13483 = n13479 & n13481 ;
  assign n13484 = n13477 | n13483 ;
  assign n31496 = ~n13484 ;
  assign n13485 = n12804 & n31496 ;
  assign n31497 = ~n12804 ;
  assign n13487 = n31497 & n13484 ;
  assign n13488 = n13485 | n13487 ;
  assign n5317 = n4246 & n5302 ;
  assign n5288 = x[109] & n5240 ;
  assign n6274 = x[110] & n6179 ;
  assign n11987 = n5288 | n6274 ;
  assign n11988 = x[111] & n5238 ;
  assign n11989 = n11987 | n11988 ;
  assign n11990 = n5317 | n11989 ;
  assign n11991 = x[23] | n11990 ;
  assign n11992 = x[23] & n11990 ;
  assign n31498 = ~n11992 ;
  assign n11993 = n11991 & n31498 ;
  assign n12568 = n12000 & n12566 ;
  assign n12574 = n12570 & n12572 ;
  assign n12575 = n12568 | n12574 ;
  assign n31499 = ~n12575 ;
  assign n12576 = n11993 & n31499 ;
  assign n31500 = ~n11993 ;
  assign n12578 = n31500 & n12575 ;
  assign n12579 = n12576 | n12578 ;
  assign n4654 = n3409 & n4632 ;
  assign n4537 = x[103] & n4514 ;
  assign n4585 = x[104] & n4572 ;
  assign n10655 = n4537 | n4585 ;
  assign n10656 = x[105] & n4504 ;
  assign n10657 = n10655 | n10656 ;
  assign n10658 = n4654 | n10657 ;
  assign n10659 = x[29] | n10658 ;
  assign n10660 = x[29] & n10658 ;
  assign n31501 = ~n10660 ;
  assign n10661 = n10659 & n31501 ;
  assign n11143 = n11132 & n11141 ;
  assign n11149 = n11145 & n11147 ;
  assign n11150 = n11143 | n11149 ;
  assign n31502 = ~n11150 ;
  assign n11151 = n10661 & n31502 ;
  assign n31503 = ~n10661 ;
  assign n11153 = n31503 & n11150 ;
  assign n11154 = n11151 | n11153 ;
  assign n4072 = n2313 & n4041 ;
  assign n3940 = x[97] & n3910 ;
  assign n4033 = x[98] & n3975 ;
  assign n9703 = n3940 | n4033 ;
  assign n9704 = x[99] & n3906 ;
  assign n9705 = n9703 | n9704 ;
  assign n9706 = n4072 | n9705 ;
  assign n31504 = ~n9706 ;
  assign n9707 = x[35] & n31504 ;
  assign n9708 = n28822 & n9706 ;
  assign n9709 = n9707 | n9708 ;
  assign n2327 = n1522 & n2321 ;
  assign n2209 = x[85] & n2179 ;
  assign n2295 = x[86] & n2244 ;
  assign n7497 = n2209 | n2295 ;
  assign n7498 = x[87] & n2175 ;
  assign n7499 = n7497 | n7498 ;
  assign n7500 = n2327 | n7499 ;
  assign n31505 = ~n7500 ;
  assign n7501 = x[47] & n31505 ;
  assign n7502 = n29621 & n7500 ;
  assign n7503 = n7501 | n7502 ;
  assign n2089 = n1457 & n2084 ;
  assign n1361 = x[76] & n1319 ;
  assign n1427 = x[77] & n1384 ;
  assign n6014 = n1361 | n1427 ;
  assign n6015 = x[78] & n1315 ;
  assign n6016 = n6014 | n6015 ;
  assign n6017 = n2089 | n6016 ;
  assign n31506 = ~n6017 ;
  assign n6018 = x[56] & n31506 ;
  assign n6019 = n30379 & n6017 ;
  assign n6020 = n6018 | n6019 ;
  assign n923 = x[70] & n900 ;
  assign n975 = x[71] & n949 ;
  assign n3697 = n923 | n975 ;
  assign n3698 = x[72] & n881 ;
  assign n3699 = n3697 | n3698 ;
  assign n3712 = n1006 & n3701 ;
  assign n3713 = n3699 | n3712 ;
  assign n31507 = ~n3713 ;
  assign n3714 = x[62] & n31507 ;
  assign n3715 = n30886 & n3713 ;
  assign n3716 = n3714 | n3715 ;
  assign n27734 = x[68] & n27215 ;
  assign n839 = x[69] & n805 ;
  assign n3694 = n27734 | n839 ;
  assign n31508 = ~n3694 ;
  assign n3695 = x[2] & n31508 ;
  assign n3717 = n27790 & n3694 ;
  assign n3718 = n3695 | n3717 ;
  assign n3719 = n3716 | n3718 ;
  assign n3720 = n3716 & n3718 ;
  assign n31509 = ~n3720 ;
  assign n4783 = n3719 & n31509 ;
  assign n4786 = x[2] & n4784 ;
  assign n4811 = n4807 & n4809 ;
  assign n4812 = n4786 | n4811 ;
  assign n4813 = n4783 | n4812 ;
  assign n4814 = n4783 & n4812 ;
  assign n31510 = ~n4814 ;
  assign n4815 = n4813 & n31510 ;
  assign n3298 = n1217 & n3289 ;
  assign n1119 = x[73] & n1079 ;
  assign n1159 = x[74] & n1144 ;
  assign n4816 = n1119 | n1159 ;
  assign n4817 = x[75] & n1075 ;
  assign n4818 = n4816 | n4817 ;
  assign n4819 = n3298 | n4818 ;
  assign n31511 = ~n4819 ;
  assign n4820 = x[59] & n31511 ;
  assign n4821 = n30638 & n4819 ;
  assign n4822 = n4820 | n4821 ;
  assign n31512 = ~n4822 ;
  assign n4823 = n4815 & n31512 ;
  assign n31513 = ~n4815 ;
  assign n5961 = n31513 & n4822 ;
  assign n5962 = n4823 | n5961 ;
  assign n5999 = n5964 & n5997 ;
  assign n6010 = n6001 & n6008 ;
  assign n6011 = n5999 | n6010 ;
  assign n6012 = n5962 | n6011 ;
  assign n6013 = n5962 & n6011 ;
  assign n31514 = ~n6013 ;
  assign n6021 = n6012 & n31514 ;
  assign n31515 = ~n6020 ;
  assign n6022 = n31515 & n6021 ;
  assign n31516 = ~n6021 ;
  assign n6371 = n6020 & n31516 ;
  assign n6372 = n6022 | n6371 ;
  assign n6538 = n6374 & n6536 ;
  assign n6549 = n6540 & n6547 ;
  assign n6550 = n6538 | n6549 ;
  assign n6551 = n6372 | n6550 ;
  assign n6552 = n6372 & n6550 ;
  assign n31517 = ~n6552 ;
  assign n6553 = n6551 & n31517 ;
  assign n1701 = n1029 & n1690 ;
  assign n1596 = x[79] & n1551 ;
  assign n1641 = x[80] & n1616 ;
  assign n6554 = n1596 | n1641 ;
  assign n6555 = x[81] & n1547 ;
  assign n6556 = n6554 | n6555 ;
  assign n6557 = n1701 | n6556 ;
  assign n31518 = ~n6557 ;
  assign n6558 = x[53] & n31518 ;
  assign n6559 = n30125 & n6557 ;
  assign n6560 = n6558 | n6559 ;
  assign n6561 = n6553 | n6560 ;
  assign n6562 = n6553 & n6560 ;
  assign n31519 = ~n6562 ;
  assign n6795 = n6561 & n31519 ;
  assign n6931 = n6921 | n6930 ;
  assign n6932 = n6795 | n6931 ;
  assign n6933 = n6795 & n6931 ;
  assign n31520 = ~n6933 ;
  assign n6934 = n6932 & n31520 ;
  assign n2025 = n1293 & n2007 ;
  assign n1919 = x[82] & n1866 ;
  assign n1986 = x[83] & n1931 ;
  assign n6935 = n1919 | n1986 ;
  assign n6936 = x[84] & n1862 ;
  assign n6937 = n6935 | n6936 ;
  assign n6938 = n2025 | n6937 ;
  assign n31521 = ~n6938 ;
  assign n6939 = x[50] & n31521 ;
  assign n6940 = n29865 & n6938 ;
  assign n6941 = n6939 | n6940 ;
  assign n31522 = ~n6941 ;
  assign n6942 = n6934 & n31522 ;
  assign n31523 = ~n6934 ;
  assign n7305 = n31523 & n6941 ;
  assign n7306 = n6942 | n7305 ;
  assign n7482 = n7308 & n7480 ;
  assign n7493 = n7484 & n7491 ;
  assign n7494 = n7482 | n7493 ;
  assign n31524 = ~n7494 ;
  assign n7495 = n7306 & n31524 ;
  assign n31525 = ~n7306 ;
  assign n7504 = n31525 & n7494 ;
  assign n7505 = n7495 | n7504 ;
  assign n31526 = ~n7503 ;
  assign n7506 = n31526 & n7505 ;
  assign n31527 = ~n7505 ;
  assign n7786 = n7503 & n31527 ;
  assign n7787 = n7506 | n7786 ;
  assign n8008 = n7789 & n8006 ;
  assign n8019 = n8010 & n8017 ;
  assign n8020 = n8008 | n8019 ;
  assign n8021 = n7787 | n8020 ;
  assign n8022 = n7787 & n8020 ;
  assign n31528 = ~n8022 ;
  assign n8023 = n8021 & n31528 ;
  assign n2655 = n1482 & n2635 ;
  assign n2545 = x[88] & n2492 ;
  assign n2609 = x[89] & n2557 ;
  assign n8024 = n2545 | n2609 ;
  assign n8025 = x[90] & n2488 ;
  assign n8026 = n8024 | n8025 ;
  assign n8027 = n2655 | n8026 ;
  assign n31529 = ~n8027 ;
  assign n8028 = x[44] & n31529 ;
  assign n8029 = n29400 & n8027 ;
  assign n8030 = n8028 | n8029 ;
  assign n31530 = ~n8030 ;
  assign n8031 = n8023 & n31530 ;
  assign n31531 = ~n8023 ;
  assign n8238 = n31531 & n8030 ;
  assign n8239 = n8031 | n8238 ;
  assign n8502 = n8241 & n8500 ;
  assign n8513 = n8504 & n8511 ;
  assign n8514 = n8502 | n8513 ;
  assign n8515 = n8239 | n8514 ;
  assign n8516 = n8239 & n8514 ;
  assign n31532 = ~n8516 ;
  assign n8517 = n8515 & n31532 ;
  assign n3177 = n1685 & n3162 ;
  assign n3036 = x[91] & n3031 ;
  assign n3142 = x[92] & n3096 ;
  assign n8518 = n3036 | n3142 ;
  assign n8519 = x[93] & n3027 ;
  assign n8520 = n8518 | n8519 ;
  assign n8521 = n3177 | n8520 ;
  assign n31533 = ~n8521 ;
  assign n8522 = x[41] & n31533 ;
  assign n8523 = n29184 & n8521 ;
  assign n8524 = n8522 | n8523 ;
  assign n31534 = ~n8524 ;
  assign n8525 = n8517 & n31534 ;
  assign n31535 = ~n8517 ;
  assign n8832 = n31535 & n8524 ;
  assign n8833 = n8525 | n8832 ;
  assign n9141 = n8835 & n9139 ;
  assign n9152 = n9143 & n9150 ;
  assign n9153 = n9141 | n9152 ;
  assign n9154 = n8833 | n9153 ;
  assign n9155 = n8833 & n9153 ;
  assign n31536 = ~n9155 ;
  assign n9156 = n9154 & n31536 ;
  assign n3589 = n2000 & n3574 ;
  assign n3501 = x[94] & n3443 ;
  assign n3510 = x[95] & n3508 ;
  assign n9157 = n3501 | n3510 ;
  assign n9158 = x[96] & n3439 ;
  assign n9159 = n9157 | n9158 ;
  assign n9160 = n3589 | n9159 ;
  assign n31537 = ~n9160 ;
  assign n9161 = x[38] & n31537 ;
  assign n9162 = n28996 & n9160 ;
  assign n9163 = n9161 | n9162 ;
  assign n31538 = ~n9163 ;
  assign n9164 = n9156 & n31538 ;
  assign n31539 = ~n9156 ;
  assign n9325 = n31539 & n9163 ;
  assign n9326 = n9164 | n9325 ;
  assign n9688 = n9328 & n9686 ;
  assign n9699 = n9690 & n9697 ;
  assign n9700 = n9688 | n9699 ;
  assign n31540 = ~n9700 ;
  assign n9701 = n9326 & n31540 ;
  assign n31541 = ~n9326 ;
  assign n9710 = n31541 & n9700 ;
  assign n9711 = n9701 | n9710 ;
  assign n31542 = ~n9709 ;
  assign n9712 = n31542 & n9711 ;
  assign n31543 = ~n9711 ;
  assign n10404 = n9709 & n31543 ;
  assign n10405 = n9712 | n10404 ;
  assign n10380 = n10376 & n10378 ;
  assign n10391 = n10387 & n10389 ;
  assign n10392 = n10380 | n10391 ;
  assign n657 = x[102] & n652 ;
  assign n10393 = x[100] & n663 ;
  assign n10394 = x[101] & n720 ;
  assign n10395 = n10393 | n10394 ;
  assign n10396 = n657 | n10395 ;
  assign n10397 = n779 & n2867 ;
  assign n10398 = n10396 | n10397 ;
  assign n10399 = n28658 & n10398 ;
  assign n31544 = ~n10398 ;
  assign n10400 = x[32] & n31544 ;
  assign n10401 = n10399 | n10400 ;
  assign n10402 = n10392 | n10401 ;
  assign n10403 = n10392 & n10401 ;
  assign n31545 = ~n10403 ;
  assign n10406 = n10402 & n31545 ;
  assign n10407 = n10405 & n10406 ;
  assign n11155 = n10405 | n10406 ;
  assign n31546 = ~n10407 ;
  assign n11156 = n31546 & n11155 ;
  assign n31547 = ~n11156 ;
  assign n11157 = n11154 & n31547 ;
  assign n31548 = ~n11154 ;
  assign n11769 = n31548 & n11156 ;
  assign n11770 = n11157 | n11769 ;
  assign n11750 = n11739 & n11748 ;
  assign n11756 = n11752 & n11754 ;
  assign n11757 = n11750 | n11756 ;
  assign n326 = x[108] & n322 ;
  assign n11758 = x[106] & n330 ;
  assign n11759 = x[107] & n390 ;
  assign n11760 = n11758 | n11759 ;
  assign n11761 = n326 | n11760 ;
  assign n11762 = n452 & n3876 ;
  assign n11763 = n11761 | n11762 ;
  assign n11764 = n28342 & n11763 ;
  assign n31549 = ~n11763 ;
  assign n11765 = x[26] & n31549 ;
  assign n11766 = n11764 | n11765 ;
  assign n31550 = ~n11766 ;
  assign n11767 = n11757 & n31550 ;
  assign n31551 = ~n11757 ;
  assign n11771 = n31551 & n11766 ;
  assign n11772 = n11767 | n11771 ;
  assign n11773 = n11770 | n11772 ;
  assign n11774 = n11770 & n11772 ;
  assign n31552 = ~n11774 ;
  assign n12580 = n11773 & n31552 ;
  assign n31553 = ~n12580 ;
  assign n12581 = n12579 & n31553 ;
  assign n31554 = ~n12579 ;
  assign n13489 = n31554 & n12580 ;
  assign n13490 = n12581 | n13489 ;
  assign n31555 = ~n13490 ;
  assign n13491 = n13488 & n31555 ;
  assign n31556 = ~n13488 ;
  assign n14293 = n31556 & n13490 ;
  assign n14294 = n13491 | n14293 ;
  assign n31557 = ~n14294 ;
  assign n14295 = n14292 & n31557 ;
  assign n31558 = ~n14292 ;
  assign n15217 = n31558 & n14294 ;
  assign n15218 = n14295 | n15217 ;
  assign n31559 = ~n15218 ;
  assign n15220 = n15216 & n31559 ;
  assign n31560 = ~n15216 ;
  assign n16276 = n31560 & n15218 ;
  assign n16277 = n15220 | n16276 ;
  assign n31561 = ~n16277 ;
  assign n17268 = n16275 & n31561 ;
  assign n31562 = ~n16275 ;
  assign n17269 = n31562 & n16277 ;
  assign n17270 = n17268 | n17269 ;
  assign n17248 = n17237 & n17246 ;
  assign n17254 = n17248 | n17253 ;
  assign n17255 = x[126] & n15244 ;
  assign n17257 = x[124] & n15246 ;
  assign n17258 = x[125] & n16288 ;
  assign n17259 = n17257 | n17258 ;
  assign n17260 = n17255 | n17259 ;
  assign n17261 = n5388 & n15308 ;
  assign n17262 = n17260 | n17261 ;
  assign n17263 = n27845 & n17262 ;
  assign n31563 = ~n17262 ;
  assign n17264 = x[8] & n31563 ;
  assign n17265 = n17263 | n17264 ;
  assign n17266 = n17254 | n17265 ;
  assign n17267 = n17254 & n17265 ;
  assign n31564 = ~n17267 ;
  assign n17271 = n17266 & n31564 ;
  assign n17272 = n17270 & n17271 ;
  assign n31565 = ~n17265 ;
  assign n18465 = n17254 & n31565 ;
  assign n31566 = ~n17254 ;
  assign n18466 = n31566 & n17265 ;
  assign n18467 = n17270 | n18466 ;
  assign n18468 = n18465 | n18467 ;
  assign n31567 = ~n17272 ;
  assign n18469 = n31567 & n18468 ;
  assign n31568 = ~n18464 ;
  assign n18470 = n31568 & n18469 ;
  assign n31569 = ~n18469 ;
  assign n18591 = n18464 & n31569 ;
  assign n18592 = n18470 | n18591 ;
  assign n31570 = ~n18592 ;
  assign n18593 = n18590 & n31570 ;
  assign n31571 = ~n18590 ;
  assign n23123 = n31571 & n18592 ;
  assign n23124 = n18593 | n23123 ;
  assign n23125 = n23122 & n23124 ;
  assign n27729 = n23122 | n23123 ;
  assign n27730 = n18593 | n27729 ;
  assign n31572 = ~n23125 ;
  assign n197 = n31572 & n27730 ;
  assign n18594 = n18590 & n18592 ;
  assign n23126 = n18594 | n23125 ;
  assign n18471 = n18464 & n18469 ;
  assign n18472 = n18463 | n18471 ;
  assign n17273 = n17267 | n17272 ;
  assign n15353 = n5629 & n15308 ;
  assign n15274 = x[125] & n15246 ;
  assign n17313 = x[126] & n16288 ;
  assign n17334 = n15274 | n17313 ;
  assign n17335 = x[127] & n15244 ;
  assign n17336 = n17334 | n17335 ;
  assign n17337 = n15353 | n17336 ;
  assign n31573 = ~n17337 ;
  assign n17338 = x[8] & n31573 ;
  assign n17339 = n27845 & n17337 ;
  assign n17340 = n17338 | n17339 ;
  assign n17341 = n17273 | n17340 ;
  assign n17342 = n17273 & n17340 ;
  assign n31574 = ~n17342 ;
  assign n17343 = n17341 & n31574 ;
  assign n12744 = n5838 & n12695 ;
  assign n12673 = x[122] & n12633 ;
  assign n14389 = x[123] & n13533 ;
  assign n15390 = n12673 | n14389 ;
  assign n15391 = x[124] & n12631 ;
  assign n15392 = n15390 | n15391 ;
  assign n15393 = n12744 | n15392 ;
  assign n31575 = ~n15393 ;
  assign n15394 = x[11] & n31575 ;
  assign n15395 = n27892 & n15393 ;
  assign n15396 = n15394 | n15395 ;
  assign n16273 = n15403 & n16271 ;
  assign n16278 = n16275 & n16277 ;
  assign n16279 = n16273 | n16278 ;
  assign n16280 = n15396 | n16279 ;
  assign n16281 = n15396 & n16279 ;
  assign n31576 = ~n16281 ;
  assign n16282 = n16280 & n31576 ;
  assign n14296 = n14292 & n14294 ;
  assign n14297 = n14291 | n14296 ;
  assign n8722 = n784 & n8706 ;
  assign n8703 = x[116] & n8645 ;
  assign n9871 = x[117] & n9278 ;
  assign n14298 = n8703 | n9871 ;
  assign n14299 = x[118] & n8643 ;
  assign n14300 = n14298 | n14299 ;
  assign n14301 = n8722 | n14300 ;
  assign n31577 = ~n14301 ;
  assign n14302 = x[17] & n31577 ;
  assign n14303 = n28039 & n14301 ;
  assign n14304 = n14302 | n14303 ;
  assign n31578 = ~n14304 ;
  assign n14305 = n14297 & n31578 ;
  assign n31579 = ~n14297 ;
  assign n14307 = n31579 & n14304 ;
  assign n14308 = n14305 | n14307 ;
  assign n5343 = n4442 & n5302 ;
  assign n5279 = x[110] & n5240 ;
  assign n6270 = x[111] & n6179 ;
  assign n11980 = n5279 | n6270 ;
  assign n11981 = x[112] & n5238 ;
  assign n11982 = n11980 | n11981 ;
  assign n11983 = n5343 | n11982 ;
  assign n11984 = x[23] | n11983 ;
  assign n11985 = x[23] & n11983 ;
  assign n31580 = ~n11985 ;
  assign n11986 = n11984 & n31580 ;
  assign n12577 = n11993 & n12575 ;
  assign n12582 = n12579 & n12580 ;
  assign n12583 = n12577 | n12582 ;
  assign n31581 = ~n12583 ;
  assign n12584 = n11986 & n31581 ;
  assign n31582 = ~n11986 ;
  assign n12586 = n31582 & n12583 ;
  assign n12587 = n12584 | n12586 ;
  assign n11768 = n11757 & n11766 ;
  assign n11775 = n11768 | n11774 ;
  assign n3640 = n452 & n3639 ;
  assign n380 = x[107] & n330 ;
  assign n403 = x[108] & n390 ;
  assign n11776 = n380 | n403 ;
  assign n11777 = x[109] & n322 ;
  assign n11778 = n11776 | n11777 ;
  assign n11779 = n3640 | n11778 ;
  assign n31583 = ~n11779 ;
  assign n11780 = x[26] & n31583 ;
  assign n11781 = n28342 & n11779 ;
  assign n11782 = n11780 | n11781 ;
  assign n11783 = n11775 | n11782 ;
  assign n11784 = n11775 & n11782 ;
  assign n31584 = ~n11784 ;
  assign n11785 = n11783 & n31584 ;
  assign n4671 = n3223 & n4632 ;
  assign n4523 = x[104] & n4514 ;
  assign n4587 = x[105] & n4572 ;
  assign n10648 = n4523 | n4587 ;
  assign n10649 = x[106] & n4504 ;
  assign n10650 = n10648 | n10649 ;
  assign n10651 = n4671 | n10650 ;
  assign n31585 = ~n10651 ;
  assign n10652 = x[29] & n31585 ;
  assign n10653 = n28483 & n10651 ;
  assign n10654 = n10652 | n10653 ;
  assign n11152 = n10661 & n11150 ;
  assign n11158 = n11154 & n11156 ;
  assign n11159 = n11152 | n11158 ;
  assign n11160 = n10654 | n11159 ;
  assign n11161 = n10654 & n11159 ;
  assign n31586 = ~n11161 ;
  assign n11162 = n11160 & n31586 ;
  assign n9702 = n9326 & n9700 ;
  assign n9713 = n9709 & n9711 ;
  assign n9714 = n9702 | n9713 ;
  assign n9165 = n9156 & n9163 ;
  assign n9166 = n9155 | n9165 ;
  assign n8526 = n8517 & n8524 ;
  assign n8527 = n8516 | n8526 ;
  assign n7496 = n7306 & n7494 ;
  assign n7507 = n7503 & n7505 ;
  assign n7508 = n7496 | n7507 ;
  assign n6943 = n6934 & n6941 ;
  assign n6944 = n6933 | n6943 ;
  assign n4824 = n4815 & n4822 ;
  assign n4825 = n4814 | n4824 ;
  assign n2758 = n1217 & n2750 ;
  assign n1112 = x[74] & n1079 ;
  assign n1190 = x[75] & n1144 ;
  assign n4772 = n1112 | n1190 ;
  assign n4773 = x[76] & n1075 ;
  assign n4774 = n4772 | n4773 ;
  assign n4775 = n2758 | n4774 ;
  assign n31587 = ~n4775 ;
  assign n4776 = x[59] & n31587 ;
  assign n4777 = n30638 & n4775 ;
  assign n4778 = n4776 | n4777 ;
  assign n3696 = x[2] & n3694 ;
  assign n3721 = n3696 | n3720 ;
  assign n27716 = x[69] & n27215 ;
  assign n829 = x[70] & n805 ;
  assign n2706 = n27716 | n829 ;
  assign n27717 = x[2] & x[5] ;
  assign n27719 = x[2] | x[5] ;
  assign n31588 = ~n27717 ;
  assign n2707 = n31588 & n27719 ;
  assign n2708 = n2706 | n2707 ;
  assign n2709 = n2706 & n2707 ;
  assign n31589 = ~n2709 ;
  assign n3722 = n2708 & n31589 ;
  assign n31590 = ~n3721 ;
  assign n3723 = n31590 & n3722 ;
  assign n31591 = ~n3722 ;
  assign n3725 = n3721 & n31591 ;
  assign n3726 = n3723 | n3725 ;
  assign n914 = x[71] & n900 ;
  assign n988 = x[72] & n949 ;
  assign n3727 = n914 | n988 ;
  assign n3728 = x[73] & n881 ;
  assign n3729 = n3727 | n3728 ;
  assign n3744 = n1006 & n3733 ;
  assign n3745 = n3729 | n3744 ;
  assign n31592 = ~n3745 ;
  assign n3746 = x[62] & n31592 ;
  assign n3747 = n30886 & n3745 ;
  assign n3748 = n3746 | n3747 ;
  assign n31593 = ~n3748 ;
  assign n3749 = n3726 & n31593 ;
  assign n31594 = ~n3726 ;
  assign n4779 = n31594 & n3748 ;
  assign n4780 = n3749 | n4779 ;
  assign n31595 = ~n4778 ;
  assign n4781 = n31595 & n4780 ;
  assign n31596 = ~n4780 ;
  assign n4826 = n4778 & n31596 ;
  assign n4827 = n4781 | n4826 ;
  assign n4828 = n4825 | n4827 ;
  assign n4829 = n4825 & n4827 ;
  assign n31597 = ~n4829 ;
  assign n5949 = n4828 & n31597 ;
  assign n1744 = n1457 & n1741 ;
  assign n1373 = x[77] & n1319 ;
  assign n1392 = x[78] & n1384 ;
  assign n5950 = n1373 | n1392 ;
  assign n5951 = x[79] & n1315 ;
  assign n5952 = n5950 | n5951 ;
  assign n5953 = n1744 | n5952 ;
  assign n31598 = ~n5953 ;
  assign n5954 = x[56] & n31598 ;
  assign n5955 = n30379 & n5953 ;
  assign n5956 = n5954 | n5955 ;
  assign n31599 = ~n5956 ;
  assign n5957 = n5949 & n31599 ;
  assign n31600 = ~n5949 ;
  assign n5959 = n31600 & n5956 ;
  assign n5960 = n5957 | n5959 ;
  assign n6023 = n6020 & n6021 ;
  assign n6024 = n6013 | n6023 ;
  assign n31601 = ~n6024 ;
  assign n6025 = n5960 & n31601 ;
  assign n31602 = ~n5960 ;
  assign n6358 = n31602 & n6024 ;
  assign n6359 = n6025 | n6358 ;
  assign n1692 = n1003 & n1690 ;
  assign n1563 = x[80] & n1551 ;
  assign n1663 = x[81] & n1616 ;
  assign n6360 = n1563 | n1663 ;
  assign n6361 = x[82] & n1547 ;
  assign n6362 = n6360 | n6361 ;
  assign n6363 = n1692 | n6362 ;
  assign n31603 = ~n6363 ;
  assign n6364 = x[53] & n31603 ;
  assign n6365 = n30125 & n6363 ;
  assign n6366 = n6364 | n6365 ;
  assign n31604 = ~n6366 ;
  assign n6367 = n6359 & n31604 ;
  assign n31605 = ~n6359 ;
  assign n6369 = n31605 & n6366 ;
  assign n6370 = n6367 | n6369 ;
  assign n6563 = n6552 | n6562 ;
  assign n31606 = ~n6563 ;
  assign n6564 = n6370 & n31606 ;
  assign n31607 = ~n6370 ;
  assign n6784 = n31607 & n6563 ;
  assign n6785 = n6564 | n6784 ;
  assign n2012 = n1239 & n2007 ;
  assign n1917 = x[83] & n1866 ;
  assign n1980 = x[84] & n1931 ;
  assign n6786 = n1917 | n1980 ;
  assign n6787 = x[85] & n1862 ;
  assign n6788 = n6786 | n6787 ;
  assign n6789 = n2012 | n6788 ;
  assign n31608 = ~n6789 ;
  assign n6790 = x[50] & n31608 ;
  assign n6791 = n29865 & n6789 ;
  assign n6792 = n6790 | n6791 ;
  assign n31609 = ~n6792 ;
  assign n6793 = n6785 & n31609 ;
  assign n31610 = ~n6785 ;
  assign n6945 = n31610 & n6792 ;
  assign n6946 = n6793 | n6945 ;
  assign n31611 = ~n6946 ;
  assign n6948 = n6944 & n31611 ;
  assign n31612 = ~n6944 ;
  assign n7294 = n31612 & n6946 ;
  assign n7295 = n6948 | n7294 ;
  assign n2331 = n1720 & n2321 ;
  assign n2220 = x[86] & n2179 ;
  assign n2293 = x[87] & n2244 ;
  assign n7296 = n2220 | n2293 ;
  assign n7297 = x[88] & n2175 ;
  assign n7298 = n7296 | n7297 ;
  assign n7299 = n2331 | n7298 ;
  assign n31613 = ~n7299 ;
  assign n7300 = x[47] & n31613 ;
  assign n7301 = n29621 & n7299 ;
  assign n7302 = n7300 | n7301 ;
  assign n7303 = n7295 | n7302 ;
  assign n7304 = n7295 & n7302 ;
  assign n31614 = ~n7304 ;
  assign n7509 = n7303 & n31614 ;
  assign n7510 = n7508 & n7509 ;
  assign n7773 = n7508 | n7509 ;
  assign n31615 = ~n7510 ;
  assign n7774 = n31615 & n7773 ;
  assign n2662 = n2046 & n2635 ;
  assign n2548 = x[89] & n2492 ;
  assign n2599 = x[90] & n2557 ;
  assign n7775 = n2548 | n2599 ;
  assign n7776 = x[91] & n2488 ;
  assign n7777 = n7775 | n7776 ;
  assign n7778 = n2662 | n7777 ;
  assign n31616 = ~n7778 ;
  assign n7779 = x[44] & n31616 ;
  assign n7780 = n29400 & n7778 ;
  assign n7781 = n7779 | n7780 ;
  assign n31617 = ~n7781 ;
  assign n7782 = n7774 & n31617 ;
  assign n31618 = ~n7774 ;
  assign n7784 = n31618 & n7781 ;
  assign n7785 = n7782 | n7784 ;
  assign n8032 = n8023 & n8030 ;
  assign n8033 = n8022 | n8032 ;
  assign n31619 = ~n8033 ;
  assign n8034 = n7785 & n31619 ;
  assign n31620 = ~n7785 ;
  assign n8228 = n31620 & n8033 ;
  assign n8229 = n8034 | n8228 ;
  assign n3181 = n2410 & n3162 ;
  assign n3086 = x[92] & n3031 ;
  assign n3123 = x[93] & n3096 ;
  assign n8230 = n3086 | n3123 ;
  assign n8231 = x[94] & n3027 ;
  assign n8232 = n8230 | n8231 ;
  assign n8233 = n3181 | n8232 ;
  assign n31621 = ~n8233 ;
  assign n8234 = x[41] & n31621 ;
  assign n8235 = n29184 & n8233 ;
  assign n8236 = n8234 | n8235 ;
  assign n8237 = n8229 & n8236 ;
  assign n8528 = n8229 | n8236 ;
  assign n31622 = ~n8237 ;
  assign n8819 = n31622 & n8528 ;
  assign n31623 = ~n8819 ;
  assign n8820 = n8527 & n31623 ;
  assign n8529 = n8527 & n8528 ;
  assign n8530 = n8237 | n8529 ;
  assign n31624 = ~n8530 ;
  assign n8821 = n8528 & n31624 ;
  assign n8822 = n8820 | n8821 ;
  assign n3579 = n2438 & n3574 ;
  assign n3497 = x[95] & n3443 ;
  assign n3564 = x[96] & n3508 ;
  assign n8823 = n3497 | n3564 ;
  assign n8824 = x[97] & n3439 ;
  assign n8825 = n8823 | n8824 ;
  assign n8826 = n3579 | n8825 ;
  assign n31625 = ~n8826 ;
  assign n8827 = x[38] & n31625 ;
  assign n8828 = n28996 & n8826 ;
  assign n8829 = n8827 | n8828 ;
  assign n31626 = ~n8829 ;
  assign n8830 = n8822 & n31626 ;
  assign n31627 = ~n8822 ;
  assign n9167 = n31627 & n8829 ;
  assign n9168 = n8830 | n9167 ;
  assign n9169 = n9166 | n9168 ;
  assign n9170 = n9166 & n9168 ;
  assign n31628 = ~n9170 ;
  assign n9315 = n9169 & n31628 ;
  assign n4064 = n2466 & n4041 ;
  assign n3958 = x[98] & n3910 ;
  assign n3989 = x[99] & n3975 ;
  assign n9316 = n3958 | n3989 ;
  assign n9317 = x[100] & n3906 ;
  assign n9318 = n9316 | n9317 ;
  assign n9319 = n4064 | n9318 ;
  assign n31629 = ~n9319 ;
  assign n9320 = x[35] & n31629 ;
  assign n9321 = n28822 & n9319 ;
  assign n9322 = n9320 | n9321 ;
  assign n9323 = n9315 | n9322 ;
  assign n9324 = n9315 & n9322 ;
  assign n31630 = ~n9324 ;
  assign n9715 = n9323 & n31630 ;
  assign n9716 = n9714 & n9715 ;
  assign n10411 = n9714 | n9715 ;
  assign n31631 = ~n9716 ;
  assign n10412 = n31631 & n10411 ;
  assign n2629 = n779 & n2626 ;
  assign n681 = x[101] & n663 ;
  assign n736 = x[102] & n720 ;
  assign n9973 = n681 | n736 ;
  assign n9974 = x[103] & n652 ;
  assign n9975 = n9973 | n9974 ;
  assign n9976 = n2629 | n9975 ;
  assign n31632 = ~n9976 ;
  assign n9977 = x[32] & n31632 ;
  assign n9978 = n28658 & n9976 ;
  assign n9979 = n9977 | n9978 ;
  assign n10408 = n10403 | n10407 ;
  assign n10409 = n9979 | n10408 ;
  assign n10410 = n9979 & n10408 ;
  assign n31633 = ~n10410 ;
  assign n10413 = n10409 & n31633 ;
  assign n10414 = n10412 & n10413 ;
  assign n11163 = n10412 | n10413 ;
  assign n31634 = ~n10414 ;
  assign n11164 = n31634 & n11163 ;
  assign n11165 = n11162 & n11164 ;
  assign n11786 = n11162 | n11164 ;
  assign n31635 = ~n11165 ;
  assign n11787 = n31635 & n11786 ;
  assign n11788 = n11785 & n11787 ;
  assign n12588 = n11785 | n11787 ;
  assign n31636 = ~n11788 ;
  assign n12589 = n31636 & n12588 ;
  assign n31637 = ~n12589 ;
  assign n12590 = n12587 & n31637 ;
  assign n31638 = ~n12587 ;
  assign n13496 = n31638 & n12589 ;
  assign n13497 = n12590 | n13496 ;
  assign n7198 = n4474 & n7162 ;
  assign n7137 = x[113] & n7100 ;
  assign n7692 = x[114] & n7647 ;
  assign n12791 = n7137 | n7692 ;
  assign n12792 = x[115] & n7098 ;
  assign n12793 = n12791 | n12792 ;
  assign n12794 = n7198 | n12793 ;
  assign n31639 = ~n12794 ;
  assign n12795 = x[20] & n31639 ;
  assign n12796 = n28114 & n12794 ;
  assign n12797 = n12795 | n12796 ;
  assign n13486 = n12804 & n13484 ;
  assign n13492 = n13488 & n13490 ;
  assign n13493 = n13486 | n13492 ;
  assign n13494 = n12797 | n13493 ;
  assign n13495 = n12797 & n13493 ;
  assign n31640 = ~n13495 ;
  assign n13498 = n13494 & n31640 ;
  assign n13499 = n13497 & n13498 ;
  assign n14309 = n13497 | n13498 ;
  assign n31641 = ~n13499 ;
  assign n14310 = n31641 & n14309 ;
  assign n14311 = n14308 | n14310 ;
  assign n14312 = n14308 & n14310 ;
  assign n31642 = ~n14312 ;
  assign n15224 = n14311 & n31642 ;
  assign n10586 = n4985 & n10542 ;
  assign n10518 = x[119] & n10481 ;
  assign n11896 = x[120] & n11232 ;
  assign n14439 = n10518 | n11896 ;
  assign n14440 = x[121] & n10479 ;
  assign n14441 = n14439 | n14440 ;
  assign n14442 = n10586 | n14441 ;
  assign n31643 = ~n14442 ;
  assign n14443 = x[14] & n31643 ;
  assign n14444 = n27956 & n14442 ;
  assign n14445 = n14443 | n14444 ;
  assign n15214 = n14452 & n15212 ;
  assign n15219 = n15216 & n15218 ;
  assign n15221 = n15214 | n15219 ;
  assign n15222 = n14445 | n15221 ;
  assign n15223 = n14445 & n15221 ;
  assign n31644 = ~n15223 ;
  assign n15225 = n15222 & n31644 ;
  assign n15226 = n15224 & n15225 ;
  assign n16283 = n15224 | n15225 ;
  assign n31645 = ~n15226 ;
  assign n16284 = n31645 & n16283 ;
  assign n16285 = n16282 | n16284 ;
  assign n16286 = n16282 & n16284 ;
  assign n31646 = ~n16286 ;
  assign n17344 = n16285 & n31646 ;
  assign n31647 = ~n17344 ;
  assign n17345 = n17343 & n31647 ;
  assign n31648 = ~n17343 ;
  assign n18473 = n31648 & n17344 ;
  assign n18474 = n17345 | n18473 ;
  assign n31649 = ~n18474 ;
  assign n18475 = n18472 & n31649 ;
  assign n31650 = ~n18472 ;
  assign n23127 = n31650 & n18474 ;
  assign n23128 = n18475 | n23127 ;
  assign n23129 = n23126 | n23128 ;
  assign n23130 = n23126 & n23128 ;
  assign n31651 = ~n23130 ;
  assign n198 = n23129 & n31651 ;
  assign n16287 = n16281 | n16286 ;
  assign n15352 = n6186 & n15308 ;
  assign n16289 = x[126] & n15246 ;
  assign n16290 = x[127] & n16288 ;
  assign n16291 = n16289 | n16290 ;
  assign n16292 = n15352 | n16291 ;
  assign n31652 = ~n16292 ;
  assign n16293 = x[8] & n31652 ;
  assign n16294 = n27845 & n16292 ;
  assign n16295 = n16293 | n16294 ;
  assign n31653 = ~n16295 ;
  assign n16296 = n16287 & n31653 ;
  assign n31654 = ~n16287 ;
  assign n16298 = n31654 & n16295 ;
  assign n16299 = n16296 | n16298 ;
  assign n12741 = n642 & n12695 ;
  assign n12679 = x[123] & n12633 ;
  assign n14390 = x[124] & n13533 ;
  assign n14432 = n12679 | n14390 ;
  assign n14433 = x[125] & n12631 ;
  assign n14434 = n14432 | n14433 ;
  assign n14435 = n12741 | n14434 ;
  assign n31655 = ~n14435 ;
  assign n14436 = x[11] & n31655 ;
  assign n14437 = n27892 & n14435 ;
  assign n14438 = n14436 | n14437 ;
  assign n15227 = n15223 | n15226 ;
  assign n15228 = n14438 | n15227 ;
  assign n15229 = n14438 & n15227 ;
  assign n31656 = ~n15229 ;
  assign n15230 = n15228 & n31656 ;
  assign n14306 = n14297 & n14304 ;
  assign n14313 = n14306 | n14312 ;
  assign n11851 = x[122] & n10479 ;
  assign n14314 = x[120] & n10481 ;
  assign n14315 = x[121] & n11232 ;
  assign n14316 = n14314 | n14315 ;
  assign n14317 = n11851 | n14316 ;
  assign n14318 = n5022 & n10542 ;
  assign n14319 = n14317 | n14318 ;
  assign n14320 = n27956 & n14319 ;
  assign n31657 = ~n14319 ;
  assign n14321 = x[14] & n31657 ;
  assign n14322 = n14320 | n14321 ;
  assign n14323 = n14313 | n14322 ;
  assign n14324 = n14313 & n14322 ;
  assign n31658 = ~n14324 ;
  assign n14325 = n14323 & n31658 ;
  assign n8746 = n5047 & n8706 ;
  assign n8684 = x[117] & n8645 ;
  assign n9857 = x[118] & n9278 ;
  assign n12784 = n8684 | n9857 ;
  assign n12785 = x[119] & n8643 ;
  assign n12786 = n12784 | n12785 ;
  assign n12787 = n8746 | n12786 ;
  assign n12788 = x[17] | n12787 ;
  assign n12789 = x[17] & n12787 ;
  assign n31659 = ~n12789 ;
  assign n12790 = n12788 & n31659 ;
  assign n13500 = n13495 | n13499 ;
  assign n31660 = ~n13500 ;
  assign n13501 = n12790 & n31660 ;
  assign n31661 = ~n12790 ;
  assign n13503 = n31661 & n13500 ;
  assign n13504 = n13501 | n13503 ;
  assign n7192 = n4702 & n7162 ;
  assign n7135 = x[114] & n7100 ;
  assign n7696 = x[115] & n7647 ;
  assign n11973 = n7135 | n7696 ;
  assign n11974 = x[116] & n7098 ;
  assign n11975 = n11973 | n11974 ;
  assign n11976 = n7192 | n11975 ;
  assign n11977 = x[20] | n11976 ;
  assign n11978 = x[20] & n11976 ;
  assign n31662 = ~n11978 ;
  assign n11979 = n11977 & n31662 ;
  assign n12585 = n11986 & n12583 ;
  assign n12591 = n12587 & n12589 ;
  assign n12592 = n12585 | n12591 ;
  assign n31663 = ~n12592 ;
  assign n12593 = n11979 & n31663 ;
  assign n31664 = ~n11979 ;
  assign n12595 = n31664 & n12592 ;
  assign n12596 = n12593 | n12595 ;
  assign n5330 = n4087 & n5302 ;
  assign n5283 = x[111] & n5240 ;
  assign n6252 = x[112] & n6179 ;
  assign n11251 = n5283 | n6252 ;
  assign n11252 = x[113] & n5238 ;
  assign n11253 = n11251 | n11252 ;
  assign n11254 = n5330 | n11253 ;
  assign n31665 = ~n11254 ;
  assign n11255 = x[23] & n31665 ;
  assign n11256 = n28221 & n11254 ;
  assign n11257 = n11255 | n11256 ;
  assign n11789 = n11784 | n11788 ;
  assign n11790 = n11257 | n11789 ;
  assign n11791 = n11257 & n11789 ;
  assign n31666 = ~n11791 ;
  assign n11792 = n11790 & n31666 ;
  assign n11166 = n11161 | n11165 ;
  assign n325 = x[110] & n322 ;
  assign n11167 = x[108] & n330 ;
  assign n11168 = x[109] & n390 ;
  assign n11169 = n11167 | n11168 ;
  assign n11170 = n325 | n11169 ;
  assign n11171 = n452 & n3615 ;
  assign n11172 = n11170 | n11171 ;
  assign n11173 = n28342 & n11172 ;
  assign n31667 = ~n11172 ;
  assign n11174 = x[26] & n31667 ;
  assign n11175 = n11173 | n11174 ;
  assign n31668 = ~n11175 ;
  assign n11176 = n11166 & n31668 ;
  assign n31669 = ~n11166 ;
  assign n11178 = n31669 & n11175 ;
  assign n11179 = n11176 | n11178 ;
  assign n4661 = n3199 & n4632 ;
  assign n4526 = x[105] & n4514 ;
  assign n4608 = x[106] & n4572 ;
  assign n9966 = n4526 | n4608 ;
  assign n9967 = x[107] & n4504 ;
  assign n9968 = n9966 | n9967 ;
  assign n9969 = n4661 | n9968 ;
  assign n9970 = x[29] | n9969 ;
  assign n9971 = x[29] & n9969 ;
  assign n31670 = ~n9971 ;
  assign n9972 = n9970 & n31670 ;
  assign n10415 = n10410 | n10414 ;
  assign n31671 = ~n10415 ;
  assign n10416 = n9972 & n31671 ;
  assign n31672 = ~n9972 ;
  assign n10418 = n31672 & n10415 ;
  assign n10419 = n10416 | n10418 ;
  assign n3002 = n779 & n3001 ;
  assign n684 = x[102] & n663 ;
  assign n733 = x[103] & n720 ;
  assign n9308 = n684 | n733 ;
  assign n9309 = x[104] & n652 ;
  assign n9310 = n9308 | n9309 ;
  assign n9311 = n3002 | n9310 ;
  assign n31673 = ~n9311 ;
  assign n9312 = x[32] & n31673 ;
  assign n9313 = n28658 & n9311 ;
  assign n9314 = n9312 | n9313 ;
  assign n9717 = n9324 | n9716 ;
  assign n9718 = n9314 | n9717 ;
  assign n9719 = n9314 & n9717 ;
  assign n31674 = ~n9719 ;
  assign n9720 = n9718 & n31674 ;
  assign n4079 = n2977 & n4041 ;
  assign n3956 = x[99] & n3910 ;
  assign n4029 = x[100] & n3975 ;
  assign n9175 = n3956 | n4029 ;
  assign n9176 = x[101] & n3906 ;
  assign n9177 = n9175 | n9176 ;
  assign n9178 = n4079 | n9177 ;
  assign n9179 = x[35] | n9178 ;
  assign n9180 = x[35] & n9178 ;
  assign n31675 = ~n9180 ;
  assign n9181 = n9179 & n31675 ;
  assign n8831 = n8822 & n8829 ;
  assign n9171 = n8831 | n9170 ;
  assign n3607 = n2841 & n3574 ;
  assign n3478 = x[96] & n3443 ;
  assign n3561 = x[97] & n3508 ;
  assign n8534 = n3478 | n3561 ;
  assign n8535 = x[98] & n3439 ;
  assign n8536 = n8534 | n8535 ;
  assign n8537 = n3607 | n8536 ;
  assign n8538 = x[38] | n8537 ;
  assign n8539 = x[38] & n8537 ;
  assign n31676 = ~n8539 ;
  assign n8540 = n8538 & n31676 ;
  assign n3724 = n3721 & n3722 ;
  assign n3750 = n3726 & n3748 ;
  assign n3751 = n3724 | n3750 ;
  assign n27714 = x[70] & n27215 ;
  assign n842 = x[71] & n805 ;
  assign n2703 = n27714 | n842 ;
  assign n2710 = n27719 & n31589 ;
  assign n31677 = ~n2703 ;
  assign n2711 = n31677 & n2710 ;
  assign n31678 = ~n2710 ;
  assign n2713 = n2703 & n31678 ;
  assign n2714 = n2711 | n2713 ;
  assign n890 = x[74] & n881 ;
  assign n2715 = x[72] & n900 ;
  assign n2716 = x[73] & n949 ;
  assign n2717 = n2715 | n2716 ;
  assign n2718 = n890 | n2717 ;
  assign n2731 = n1006 & n2722 ;
  assign n2732 = n2718 | n2731 ;
  assign n2733 = n30886 & n2732 ;
  assign n31679 = ~n2732 ;
  assign n2734 = x[62] & n31679 ;
  assign n2735 = n2733 | n2734 ;
  assign n31680 = ~n2735 ;
  assign n2736 = n2714 & n31680 ;
  assign n31681 = ~n2714 ;
  assign n3752 = n31681 & n2735 ;
  assign n3753 = n2736 | n3752 ;
  assign n31682 = ~n3751 ;
  assign n3754 = n31682 & n3753 ;
  assign n31683 = ~n3753 ;
  assign n3756 = n3751 & n31683 ;
  assign n3757 = n3754 | n3756 ;
  assign n1780 = n1217 & n1775 ;
  assign n1108 = x[75] & n1079 ;
  assign n1201 = x[76] & n1144 ;
  assign n3758 = n1108 | n1201 ;
  assign n3759 = x[77] & n1075 ;
  assign n3760 = n3758 | n3759 ;
  assign n3761 = n1780 | n3760 ;
  assign n31684 = ~n3761 ;
  assign n3762 = x[59] & n31684 ;
  assign n3763 = n30638 & n3761 ;
  assign n3764 = n3762 | n3763 ;
  assign n31685 = ~n3764 ;
  assign n3765 = n3757 & n31685 ;
  assign n31686 = ~n3757 ;
  assign n4770 = n31686 & n3764 ;
  assign n4771 = n3765 | n4770 ;
  assign n4782 = n4778 & n4780 ;
  assign n4830 = n4782 | n4829 ;
  assign n4831 = n4771 | n4830 ;
  assign n4832 = n4771 & n4830 ;
  assign n31687 = ~n4832 ;
  assign n4833 = n4831 & n31687 ;
  assign n1464 = n1270 & n1457 ;
  assign n1355 = x[78] & n1319 ;
  assign n1390 = x[79] & n1384 ;
  assign n4834 = n1355 | n1390 ;
  assign n4835 = x[80] & n1315 ;
  assign n4836 = n4834 | n4835 ;
  assign n4837 = n1464 | n4836 ;
  assign n31688 = ~n4837 ;
  assign n4838 = x[56] & n31688 ;
  assign n4839 = n30379 & n4837 ;
  assign n4840 = n4838 | n4839 ;
  assign n31689 = ~n4840 ;
  assign n4841 = n4833 & n31689 ;
  assign n31690 = ~n4833 ;
  assign n5947 = n31690 & n4840 ;
  assign n5948 = n4841 | n5947 ;
  assign n5958 = n5949 & n5956 ;
  assign n6026 = n5960 & n6024 ;
  assign n6027 = n5958 | n6026 ;
  assign n6028 = n5948 | n6027 ;
  assign n6029 = n5948 & n6027 ;
  assign n31691 = ~n6029 ;
  assign n6030 = n6028 & n31691 ;
  assign n1699 = n1057 & n1690 ;
  assign n1604 = x[81] & n1551 ;
  assign n1671 = x[82] & n1616 ;
  assign n6031 = n1604 | n1671 ;
  assign n6032 = x[83] & n1547 ;
  assign n6033 = n6031 | n6032 ;
  assign n6034 = n1699 | n6033 ;
  assign n31692 = ~n6034 ;
  assign n6035 = x[53] & n31692 ;
  assign n6036 = n30125 & n6034 ;
  assign n6037 = n6035 | n6036 ;
  assign n31693 = ~n6037 ;
  assign n6038 = n6030 & n31693 ;
  assign n31694 = ~n6030 ;
  assign n6356 = n31694 & n6037 ;
  assign n6357 = n6038 | n6356 ;
  assign n6368 = n6359 & n6366 ;
  assign n6565 = n6370 & n6563 ;
  assign n6566 = n6368 | n6565 ;
  assign n6567 = n6357 | n6566 ;
  assign n6568 = n6357 & n6566 ;
  assign n31695 = ~n6568 ;
  assign n6569 = n6567 & n31695 ;
  assign n2024 = n1213 & n2007 ;
  assign n1910 = x[84] & n1866 ;
  assign n1950 = x[85] & n1931 ;
  assign n6570 = n1910 | n1950 ;
  assign n6571 = x[86] & n1862 ;
  assign n6572 = n6570 | n6571 ;
  assign n6573 = n2024 | n6572 ;
  assign n31696 = ~n6573 ;
  assign n6574 = x[50] & n31696 ;
  assign n6575 = n29865 & n6573 ;
  assign n6576 = n6574 | n6575 ;
  assign n31697 = ~n6576 ;
  assign n6577 = n6569 & n31697 ;
  assign n31698 = ~n6569 ;
  assign n6782 = n31698 & n6576 ;
  assign n6783 = n6577 | n6782 ;
  assign n6794 = n6785 & n6792 ;
  assign n6947 = n6944 & n6946 ;
  assign n6949 = n6794 | n6947 ;
  assign n31699 = ~n6949 ;
  assign n6950 = n6783 & n31699 ;
  assign n31700 = ~n6783 ;
  assign n6952 = n31700 & n6949 ;
  assign n6953 = n6950 | n6952 ;
  assign n2328 = n1453 & n2321 ;
  assign n2213 = x[87] & n2179 ;
  assign n2280 = x[88] & n2244 ;
  assign n6954 = n2213 | n2280 ;
  assign n6955 = x[89] & n2175 ;
  assign n6956 = n6954 | n6955 ;
  assign n6957 = n2328 | n6956 ;
  assign n31701 = ~n6957 ;
  assign n6958 = x[47] & n31701 ;
  assign n6959 = n29621 & n6957 ;
  assign n6960 = n6958 | n6959 ;
  assign n31702 = ~n6960 ;
  assign n6961 = n6953 & n31702 ;
  assign n31703 = ~n6953 ;
  assign n7292 = n31703 & n6960 ;
  assign n7293 = n6961 | n7292 ;
  assign n7511 = n7304 | n7510 ;
  assign n31704 = ~n7511 ;
  assign n7512 = n7293 & n31704 ;
  assign n31705 = ~n7293 ;
  assign n7514 = n31705 & n7511 ;
  assign n7515 = n7512 | n7514 ;
  assign n2656 = n1841 & n2635 ;
  assign n2536 = x[90] & n2492 ;
  assign n2604 = x[91] & n2557 ;
  assign n7516 = n2536 | n2604 ;
  assign n7517 = x[92] & n2488 ;
  assign n7518 = n7516 | n7517 ;
  assign n7519 = n2656 | n7518 ;
  assign n31706 = ~n7519 ;
  assign n7520 = x[44] & n31706 ;
  assign n7521 = n29400 & n7519 ;
  assign n7522 = n7520 | n7521 ;
  assign n31707 = ~n7522 ;
  assign n7523 = n7515 & n31707 ;
  assign n31708 = ~n7515 ;
  assign n7771 = n31708 & n7522 ;
  assign n7772 = n7523 | n7771 ;
  assign n7783 = n7774 & n7781 ;
  assign n8035 = n7785 & n8033 ;
  assign n8036 = n7783 | n8035 ;
  assign n31709 = ~n8036 ;
  assign n8037 = n7772 & n31709 ;
  assign n31710 = ~n7772 ;
  assign n8039 = n31710 & n8036 ;
  assign n8040 = n8037 | n8039 ;
  assign n3194 = n2152 & n3162 ;
  assign n3066 = x[93] & n3031 ;
  assign n3147 = x[94] & n3096 ;
  assign n8041 = n3066 | n3147 ;
  assign n8042 = x[95] & n3027 ;
  assign n8043 = n8041 | n8042 ;
  assign n8044 = n3194 | n8043 ;
  assign n31711 = ~n8044 ;
  assign n8045 = x[41] & n31711 ;
  assign n8046 = n29184 & n8044 ;
  assign n8047 = n8045 | n8046 ;
  assign n31712 = ~n8047 ;
  assign n8048 = n8040 & n31712 ;
  assign n31713 = ~n8040 ;
  assign n8531 = n31713 & n8047 ;
  assign n8532 = n8048 | n8531 ;
  assign n8533 = n8530 & n8532 ;
  assign n8541 = n8530 | n8532 ;
  assign n31714 = ~n8533 ;
  assign n8542 = n31714 & n8541 ;
  assign n8543 = n8540 & n8542 ;
  assign n9172 = n8540 | n8542 ;
  assign n31715 = ~n8543 ;
  assign n9173 = n31715 & n9172 ;
  assign n9174 = n9171 & n9173 ;
  assign n9182 = n9171 | n9173 ;
  assign n31716 = ~n9174 ;
  assign n9183 = n31716 & n9182 ;
  assign n9184 = n9181 & n9183 ;
  assign n9721 = n9181 | n9183 ;
  assign n31717 = ~n9184 ;
  assign n9722 = n31717 & n9721 ;
  assign n31718 = ~n9722 ;
  assign n9723 = n9720 & n31718 ;
  assign n31719 = ~n9720 ;
  assign n10420 = n31719 & n9722 ;
  assign n10421 = n9723 | n10420 ;
  assign n31720 = ~n10421 ;
  assign n10423 = n10419 & n31720 ;
  assign n31721 = ~n10419 ;
  assign n11180 = n31721 & n10421 ;
  assign n11181 = n10423 | n11180 ;
  assign n31722 = ~n11181 ;
  assign n11182 = n11179 & n31722 ;
  assign n31723 = ~n11179 ;
  assign n11793 = n31723 & n11181 ;
  assign n11794 = n11182 | n11793 ;
  assign n31724 = ~n11794 ;
  assign n11795 = n11792 & n31724 ;
  assign n31725 = ~n11792 ;
  assign n12597 = n31725 & n11794 ;
  assign n12598 = n11795 | n12597 ;
  assign n31726 = ~n12598 ;
  assign n12599 = n12596 & n31726 ;
  assign n31727 = ~n12596 ;
  assign n13505 = n31727 & n12598 ;
  assign n13506 = n12599 | n13505 ;
  assign n13507 = n13504 & n13506 ;
  assign n14326 = n13504 | n13506 ;
  assign n31728 = ~n13507 ;
  assign n14327 = n31728 & n14326 ;
  assign n31729 = ~n14327 ;
  assign n15231 = n14325 & n31729 ;
  assign n15232 = n31728 & n14325 ;
  assign n31730 = ~n15232 ;
  assign n15233 = n14326 & n31730 ;
  assign n15234 = n31728 & n15233 ;
  assign n15235 = n15231 | n15234 ;
  assign n15236 = n15230 & n15235 ;
  assign n16300 = n15230 | n15235 ;
  assign n31731 = ~n15236 ;
  assign n16307 = n31731 & n16300 ;
  assign n31732 = ~n16307 ;
  assign n16308 = n16299 & n31732 ;
  assign n16309 = n31731 & n16299 ;
  assign n31733 = ~n16309 ;
  assign n16310 = n16300 & n31733 ;
  assign n16311 = n31731 & n16310 ;
  assign n16312 = n16308 | n16311 ;
  assign n17346 = n17343 & n17344 ;
  assign n17347 = n17342 | n17346 ;
  assign n31734 = ~n17347 ;
  assign n17348 = n16312 & n31734 ;
  assign n31735 = ~n16312 ;
  assign n17350 = n31735 & n17347 ;
  assign n17351 = n17348 | n17350 ;
  assign n18476 = n18472 & n18474 ;
  assign n23131 = n18476 | n23130 ;
  assign n23132 = n17351 & n23131 ;
  assign n27733 = n17351 | n23131 ;
  assign n31736 = ~n23132 ;
  assign n199 = n31736 & n27733 ;
  assign n17349 = n16312 & n17347 ;
  assign n23133 = n17349 | n23132 ;
  assign n16297 = n16287 & n16295 ;
  assign n16301 = n16299 & n16300 ;
  assign n16302 = n31731 & n16301 ;
  assign n16303 = n16297 | n16302 ;
  assign n15237 = n15229 | n15236 ;
  assign n15288 = x[127] & n15246 ;
  assign n15354 = n5360 & n15308 ;
  assign n15372 = n15288 | n15354 ;
  assign n31737 = ~n15372 ;
  assign n15373 = x[8] & n31737 ;
  assign n15374 = n27845 & n15372 ;
  assign n15375 = n15373 | n15374 ;
  assign n31738 = ~n15375 ;
  assign n15376 = n15237 & n31738 ;
  assign n31739 = ~n15237 ;
  assign n15378 = n31739 & n15375 ;
  assign n15379 = n15376 | n15378 ;
  assign n8754 = n4678 & n8706 ;
  assign n8686 = x[118] & n8645 ;
  assign n9866 = x[119] & n9278 ;
  assign n11966 = n8686 | n9866 ;
  assign n11967 = x[120] & n8643 ;
  assign n11968 = n11966 | n11967 ;
  assign n11969 = n8754 | n11968 ;
  assign n11970 = x[17] | n11969 ;
  assign n11971 = x[17] & n11969 ;
  assign n31740 = ~n11971 ;
  assign n11972 = n11970 & n31740 ;
  assign n12594 = n11979 & n12592 ;
  assign n12600 = n12596 & n12598 ;
  assign n12601 = n12594 | n12600 ;
  assign n31741 = ~n12601 ;
  assign n12602 = n11972 & n31741 ;
  assign n31742 = ~n11972 ;
  assign n12604 = n31742 & n12601 ;
  assign n12605 = n12602 | n12604 ;
  assign n5347 = n4276 & n5302 ;
  assign n5249 = x[112] & n5240 ;
  assign n6276 = x[113] & n6179 ;
  assign n10641 = n5249 | n6276 ;
  assign n10642 = x[114] & n5238 ;
  assign n10643 = n10641 | n10642 ;
  assign n10644 = n5347 | n10643 ;
  assign n10645 = x[23] | n10644 ;
  assign n10646 = x[23] & n10644 ;
  assign n31743 = ~n10646 ;
  assign n10647 = n10645 & n31743 ;
  assign n11177 = n11166 & n11175 ;
  assign n11183 = n11179 & n11181 ;
  assign n11184 = n11177 | n11183 ;
  assign n31744 = ~n11184 ;
  assign n11185 = n10647 & n31744 ;
  assign n31745 = ~n10647 ;
  assign n11187 = n31745 & n11184 ;
  assign n11188 = n11185 | n11187 ;
  assign n4247 = n452 & n4246 ;
  assign n385 = x[109] & n330 ;
  assign n394 = x[110] & n390 ;
  assign n9959 = n385 | n394 ;
  assign n9960 = x[111] & n322 ;
  assign n9961 = n9959 | n9960 ;
  assign n9962 = n4247 | n9961 ;
  assign n31746 = ~n9962 ;
  assign n9963 = x[26] & n31746 ;
  assign n9964 = n28342 & n9962 ;
  assign n9965 = n9963 | n9964 ;
  assign n10417 = n9972 & n10415 ;
  assign n10422 = n10419 & n10421 ;
  assign n10424 = n10417 | n10422 ;
  assign n31747 = ~n10424 ;
  assign n10425 = n9965 & n31747 ;
  assign n31748 = ~n9965 ;
  assign n10427 = n31748 & n10424 ;
  assign n10428 = n10425 | n10427 ;
  assign n3413 = n779 & n3409 ;
  assign n683 = x[103] & n663 ;
  assign n742 = x[104] & n720 ;
  assign n8812 = n683 | n742 ;
  assign n8813 = x[105] & n652 ;
  assign n8814 = n8812 | n8813 ;
  assign n8815 = n3413 | n8814 ;
  assign n31749 = ~n8815 ;
  assign n8816 = x[32] & n31749 ;
  assign n8817 = n28658 & n8815 ;
  assign n8818 = n8816 | n8817 ;
  assign n9185 = n9174 | n9184 ;
  assign n31750 = ~n9185 ;
  assign n9186 = n8818 & n31750 ;
  assign n31751 = ~n8818 ;
  assign n9188 = n31751 & n9185 ;
  assign n9189 = n9186 | n9188 ;
  assign n3606 = n2313 & n3574 ;
  assign n3496 = x[97] & n3443 ;
  assign n3559 = x[98] & n3508 ;
  assign n8053 = n3496 | n3559 ;
  assign n8054 = x[99] & n3439 ;
  assign n8055 = n8053 | n8054 ;
  assign n8056 = n3606 | n8055 ;
  assign n31752 = ~n8056 ;
  assign n8057 = x[38] & n31752 ;
  assign n8058 = n28996 & n8056 ;
  assign n8059 = n8057 | n8058 ;
  assign n2338 = n1482 & n2321 ;
  assign n2227 = x[88] & n2179 ;
  assign n2292 = x[89] & n2244 ;
  assign n6585 = n2227 | n2292 ;
  assign n6586 = x[90] & n2175 ;
  assign n6587 = n6585 | n6586 ;
  assign n6588 = n2338 | n6587 ;
  assign n31753 = ~n6588 ;
  assign n6589 = x[47] & n31753 ;
  assign n6590 = n29621 & n6588 ;
  assign n6591 = n6589 | n6590 ;
  assign n6578 = n6569 & n6576 ;
  assign n6579 = n6568 | n6578 ;
  assign n2023 = n1522 & n2007 ;
  assign n1922 = x[85] & n1866 ;
  assign n1970 = x[86] & n1931 ;
  assign n6044 = n1922 | n1970 ;
  assign n6045 = x[87] & n1862 ;
  assign n6046 = n6044 | n6045 ;
  assign n6047 = n2023 | n6046 ;
  assign n6048 = x[50] | n6047 ;
  assign n6049 = x[50] & n6047 ;
  assign n31754 = ~n6049 ;
  assign n6050 = n6048 & n31754 ;
  assign n6039 = n6030 & n6037 ;
  assign n6040 = n6029 | n6039 ;
  assign n3755 = n3751 & n3753 ;
  assign n3766 = n3757 & n3764 ;
  assign n3767 = n3755 | n3766 ;
  assign n2712 = n2703 | n2710 ;
  assign n2737 = n2714 & n2735 ;
  assign n31755 = ~n2737 ;
  assign n2738 = n2712 & n31755 ;
  assign n27694 = x[71] & n27215 ;
  assign n864 = x[72] & n805 ;
  assign n1759 = n27694 | n864 ;
  assign n31756 = ~n1759 ;
  assign n2704 = n31756 & n2703 ;
  assign n2705 = n1759 & n31677 ;
  assign n3279 = n2704 | n2705 ;
  assign n31757 = ~n2738 ;
  assign n3280 = n31757 & n3279 ;
  assign n2739 = n2705 | n2738 ;
  assign n31758 = ~n2704 ;
  assign n2740 = n31758 & n2739 ;
  assign n31759 = ~n2705 ;
  assign n3281 = n31759 & n2740 ;
  assign n3282 = n3280 | n3281 ;
  assign n936 = x[73] & n900 ;
  assign n978 = x[74] & n949 ;
  assign n3283 = n936 | n978 ;
  assign n3284 = x[75] & n881 ;
  assign n3285 = n3283 | n3284 ;
  assign n3299 = n1006 & n3289 ;
  assign n3300 = n3285 | n3299 ;
  assign n31760 = ~n3300 ;
  assign n3301 = x[62] & n31760 ;
  assign n3302 = n30886 & n3300 ;
  assign n3303 = n3301 | n3302 ;
  assign n31761 = ~n3303 ;
  assign n3304 = n3282 & n31761 ;
  assign n31762 = ~n3282 ;
  assign n3305 = n31762 & n3303 ;
  assign n3306 = n3304 | n3305 ;
  assign n2090 = n1217 & n2084 ;
  assign n1117 = x[76] & n1079 ;
  assign n1149 = x[77] & n1144 ;
  assign n3307 = n1117 | n1149 ;
  assign n3308 = x[78] & n1075 ;
  assign n3309 = n3307 | n3308 ;
  assign n3310 = n2090 | n3309 ;
  assign n31763 = ~n3310 ;
  assign n3311 = x[59] & n31763 ;
  assign n3312 = n30638 & n3310 ;
  assign n3313 = n3311 | n3312 ;
  assign n3314 = n3306 | n3313 ;
  assign n3316 = n3306 & n3313 ;
  assign n31764 = ~n3316 ;
  assign n3768 = n3314 & n31764 ;
  assign n3769 = n3767 & n3768 ;
  assign n3770 = n3767 | n3768 ;
  assign n31765 = ~n3769 ;
  assign n3771 = n31765 & n3770 ;
  assign n1459 = n1029 & n1457 ;
  assign n1357 = x[79] & n1319 ;
  assign n1411 = x[80] & n1384 ;
  assign n3772 = n1357 | n1411 ;
  assign n3773 = x[81] & n1315 ;
  assign n3774 = n3772 | n3773 ;
  assign n3775 = n1459 | n3774 ;
  assign n31766 = ~n3775 ;
  assign n3776 = x[56] & n31766 ;
  assign n3777 = n30379 & n3775 ;
  assign n3778 = n3776 | n3777 ;
  assign n31767 = ~n3778 ;
  assign n3779 = n3771 & n31767 ;
  assign n31768 = ~n3771 ;
  assign n4768 = n31768 & n3778 ;
  assign n4769 = n3779 | n4768 ;
  assign n4842 = n4833 & n4840 ;
  assign n4843 = n4832 | n4842 ;
  assign n4844 = n4769 | n4843 ;
  assign n4845 = n4769 & n4843 ;
  assign n31769 = ~n4845 ;
  assign n4846 = n4844 & n31769 ;
  assign n1700 = n1293 & n1690 ;
  assign n1598 = x[82] & n1551 ;
  assign n1667 = x[83] & n1616 ;
  assign n4847 = n1598 | n1667 ;
  assign n4848 = x[84] & n1547 ;
  assign n4849 = n4847 | n4848 ;
  assign n4850 = n1700 | n4849 ;
  assign n31770 = ~n4850 ;
  assign n4851 = x[53] & n31770 ;
  assign n4852 = n30125 & n4850 ;
  assign n4853 = n4851 | n4852 ;
  assign n31771 = ~n4853 ;
  assign n4854 = n4846 & n31771 ;
  assign n31772 = ~n4846 ;
  assign n6041 = n31772 & n4853 ;
  assign n6042 = n4854 | n6041 ;
  assign n31773 = ~n6042 ;
  assign n6051 = n6040 & n31773 ;
  assign n31774 = ~n6040 ;
  assign n6052 = n31774 & n6042 ;
  assign n6053 = n6051 | n6052 ;
  assign n6054 = n6050 & n6053 ;
  assign n6580 = n6050 | n6052 ;
  assign n6581 = n6051 | n6580 ;
  assign n31775 = ~n6054 ;
  assign n6582 = n31775 & n6581 ;
  assign n6583 = n6579 | n6582 ;
  assign n6584 = n6579 & n6582 ;
  assign n31776 = ~n6584 ;
  assign n6592 = n6583 & n31776 ;
  assign n31777 = ~n6591 ;
  assign n6594 = n31777 & n6592 ;
  assign n31778 = ~n6592 ;
  assign n6780 = n6591 & n31778 ;
  assign n6781 = n6594 | n6780 ;
  assign n6951 = n6783 & n6949 ;
  assign n6962 = n6953 & n6960 ;
  assign n6963 = n6951 | n6962 ;
  assign n6964 = n6781 | n6963 ;
  assign n6965 = n6781 & n6963 ;
  assign n31779 = ~n6965 ;
  assign n6966 = n6964 & n31779 ;
  assign n2653 = n1685 & n2635 ;
  assign n2547 = x[91] & n2492 ;
  assign n2591 = x[92] & n2557 ;
  assign n6967 = n2547 | n2591 ;
  assign n6968 = x[93] & n2488 ;
  assign n6969 = n6967 | n6968 ;
  assign n6970 = n2653 | n6969 ;
  assign n31780 = ~n6970 ;
  assign n6971 = x[44] & n31780 ;
  assign n6972 = n29400 & n6970 ;
  assign n6973 = n6971 | n6972 ;
  assign n31781 = ~n6973 ;
  assign n6974 = n6966 & n31781 ;
  assign n31782 = ~n6966 ;
  assign n7290 = n31782 & n6973 ;
  assign n7291 = n6974 | n7290 ;
  assign n7513 = n7293 & n7511 ;
  assign n7524 = n7515 & n7522 ;
  assign n7525 = n7513 | n7524 ;
  assign n7526 = n7291 | n7525 ;
  assign n7527 = n7291 & n7525 ;
  assign n31783 = ~n7527 ;
  assign n7528 = n7526 & n31783 ;
  assign n3174 = n2000 & n3162 ;
  assign n3078 = x[94] & n3031 ;
  assign n3134 = x[95] & n3096 ;
  assign n7529 = n3078 | n3134 ;
  assign n7530 = x[96] & n3027 ;
  assign n7531 = n7529 | n7530 ;
  assign n7532 = n3174 | n7531 ;
  assign n31784 = ~n7532 ;
  assign n7533 = x[41] & n31784 ;
  assign n7534 = n29184 & n7532 ;
  assign n7535 = n7533 | n7534 ;
  assign n31785 = ~n7535 ;
  assign n7536 = n7528 & n31785 ;
  assign n31786 = ~n7528 ;
  assign n7769 = n31786 & n7535 ;
  assign n7770 = n7536 | n7769 ;
  assign n8038 = n7772 & n8036 ;
  assign n8049 = n8040 & n8047 ;
  assign n8050 = n8038 | n8049 ;
  assign n31787 = ~n8050 ;
  assign n8051 = n7770 & n31787 ;
  assign n31788 = ~n7770 ;
  assign n8060 = n31788 & n8050 ;
  assign n8061 = n8051 | n8060 ;
  assign n31789 = ~n8059 ;
  assign n8063 = n31789 & n8061 ;
  assign n31790 = ~n8061 ;
  assign n8226 = n8059 & n31790 ;
  assign n8227 = n8063 | n8226 ;
  assign n8544 = n8533 | n8543 ;
  assign n8545 = n8227 | n8544 ;
  assign n8546 = n8227 & n8544 ;
  assign n31791 = ~n8546 ;
  assign n8547 = n8545 & n31791 ;
  assign n4070 = n2867 & n4041 ;
  assign n3953 = x[100] & n3910 ;
  assign n3991 = x[101] & n3975 ;
  assign n8548 = n3953 | n3991 ;
  assign n8549 = x[102] & n3906 ;
  assign n8550 = n8548 | n8549 ;
  assign n8551 = n4070 | n8550 ;
  assign n31792 = ~n8551 ;
  assign n8552 = x[35] & n31792 ;
  assign n8553 = n28822 & n8551 ;
  assign n8554 = n8552 | n8553 ;
  assign n8555 = n8547 & n8554 ;
  assign n9190 = n8547 | n8554 ;
  assign n9191 = n9189 & n9190 ;
  assign n31793 = ~n8555 ;
  assign n9192 = n31793 & n9191 ;
  assign n31794 = ~n9192 ;
  assign n9737 = n9189 & n31794 ;
  assign n9738 = n9190 & n31794 ;
  assign n9739 = n31793 & n9738 ;
  assign n9740 = n9737 | n9739 ;
  assign n9724 = n9720 & n9722 ;
  assign n9725 = n9719 | n9724 ;
  assign n4509 = x[108] & n4504 ;
  assign n9726 = x[106] & n4514 ;
  assign n9727 = x[107] & n4572 ;
  assign n9728 = n9726 | n9727 ;
  assign n9729 = n4509 | n9728 ;
  assign n9730 = n3876 & n4632 ;
  assign n9731 = n9729 | n9730 ;
  assign n9732 = n28483 & n9731 ;
  assign n31795 = ~n9731 ;
  assign n9733 = x[29] & n31795 ;
  assign n9734 = n9732 | n9733 ;
  assign n9735 = n9725 | n9734 ;
  assign n9736 = n9725 & n9734 ;
  assign n31796 = ~n9736 ;
  assign n9741 = n9735 & n31796 ;
  assign n9742 = n9740 | n9741 ;
  assign n9743 = n9740 & n9741 ;
  assign n31797 = ~n9743 ;
  assign n10429 = n9742 & n31797 ;
  assign n10430 = n10428 | n10429 ;
  assign n10431 = n10428 & n10429 ;
  assign n31798 = ~n10431 ;
  assign n11189 = n10430 & n31798 ;
  assign n31799 = ~n11189 ;
  assign n11190 = n11188 & n31799 ;
  assign n31800 = ~n11188 ;
  assign n11809 = n31800 & n11189 ;
  assign n11810 = n11190 | n11809 ;
  assign n11796 = n11792 & n11794 ;
  assign n11797 = n11791 | n11796 ;
  assign n7670 = x[117] & n7098 ;
  assign n11798 = x[115] & n7100 ;
  assign n11799 = x[116] & n7647 ;
  assign n11800 = n11798 | n11799 ;
  assign n11801 = n7670 | n11800 ;
  assign n11802 = n797 & n7162 ;
  assign n11803 = n11801 | n11802 ;
  assign n11804 = n28114 & n11803 ;
  assign n31801 = ~n11803 ;
  assign n11805 = x[20] & n31801 ;
  assign n11806 = n11804 | n11805 ;
  assign n31802 = ~n11806 ;
  assign n11807 = n11797 & n31802 ;
  assign n31803 = ~n11797 ;
  assign n11811 = n31803 & n11806 ;
  assign n11812 = n11807 | n11811 ;
  assign n31804 = ~n11812 ;
  assign n11813 = n11810 & n31804 ;
  assign n31805 = ~n11810 ;
  assign n12606 = n31805 & n11812 ;
  assign n12607 = n11813 | n12606 ;
  assign n31806 = ~n12607 ;
  assign n12608 = n12605 & n31806 ;
  assign n31807 = ~n12605 ;
  assign n13511 = n31807 & n12607 ;
  assign n13512 = n12608 | n13511 ;
  assign n10579 = n5417 & n10542 ;
  assign n10519 = x[121] & n10481 ;
  assign n11904 = x[122] & n11232 ;
  assign n12777 = n10519 | n11904 ;
  assign n12778 = x[123] & n10479 ;
  assign n12779 = n12777 | n12778 ;
  assign n12780 = n10579 | n12779 ;
  assign n31808 = ~n12780 ;
  assign n12781 = x[14] & n31808 ;
  assign n12782 = n27956 & n12780 ;
  assign n12783 = n12781 | n12782 ;
  assign n13502 = n12790 & n13500 ;
  assign n13508 = n13502 | n13507 ;
  assign n31809 = ~n13508 ;
  assign n13509 = n12783 & n31809 ;
  assign n31810 = ~n12783 ;
  assign n13513 = n31810 & n13508 ;
  assign n13514 = n13509 | n13513 ;
  assign n13515 = n13512 | n13514 ;
  assign n13516 = n13512 & n13514 ;
  assign n31811 = ~n13516 ;
  assign n14344 = n13515 & n31811 ;
  assign n14328 = n14325 & n14326 ;
  assign n14329 = n31728 & n14328 ;
  assign n14330 = n14324 | n14329 ;
  assign n14331 = x[126] & n12631 ;
  assign n14333 = x[124] & n12633 ;
  assign n14334 = x[125] & n13533 ;
  assign n14335 = n14333 | n14334 ;
  assign n14336 = n14331 | n14335 ;
  assign n14337 = n5388 & n12695 ;
  assign n14338 = n14336 | n14337 ;
  assign n14339 = n27892 & n14338 ;
  assign n31812 = ~n14338 ;
  assign n14340 = x[11] & n31812 ;
  assign n14341 = n14339 | n14340 ;
  assign n14343 = n14330 & n14341 ;
  assign n14345 = n14330 | n14341 ;
  assign n31813 = ~n14343 ;
  assign n14347 = n31813 & n14345 ;
  assign n14348 = n14344 & n14347 ;
  assign n31814 = ~n14341 ;
  assign n14342 = n14330 & n31814 ;
  assign n31815 = ~n14330 ;
  assign n14346 = n31815 & n14341 ;
  assign n15380 = n14344 | n14346 ;
  assign n15381 = n14342 | n15380 ;
  assign n31816 = ~n14348 ;
  assign n15382 = n31816 & n15381 ;
  assign n31817 = ~n15379 ;
  assign n15383 = n31817 & n15382 ;
  assign n31818 = ~n15382 ;
  assign n16304 = n15379 & n31818 ;
  assign n16305 = n15383 | n16304 ;
  assign n31819 = ~n16305 ;
  assign n23134 = n16303 & n31819 ;
  assign n31820 = ~n16303 ;
  assign n23135 = n31820 & n16305 ;
  assign n23136 = n23134 | n23135 ;
  assign n23137 = n23133 & n23136 ;
  assign n27735 = n23133 | n23135 ;
  assign n27736 = n23134 | n27735 ;
  assign n31821 = ~n23137 ;
  assign n200 = n31821 & n27736 ;
  assign n16306 = n16303 & n16305 ;
  assign n23138 = n16306 | n23137 ;
  assign n15377 = n15237 & n15375 ;
  assign n15384 = n15379 & n15382 ;
  assign n15385 = n15377 | n15384 ;
  assign n14349 = n14343 | n14348 ;
  assign n12743 = n5629 & n12695 ;
  assign n12667 = x[125] & n12633 ;
  assign n14380 = x[126] & n13533 ;
  assign n14410 = n12667 | n14380 ;
  assign n14411 = x[127] & n12631 ;
  assign n14412 = n14410 | n14411 ;
  assign n14413 = n12743 | n14412 ;
  assign n31822 = ~n14413 ;
  assign n14414 = x[11] & n31822 ;
  assign n14415 = n27892 & n14413 ;
  assign n14416 = n14414 | n14415 ;
  assign n14417 = n14349 | n14416 ;
  assign n14418 = n14349 & n14416 ;
  assign n31823 = ~n14418 ;
  assign n14419 = n14417 & n31823 ;
  assign n13510 = n12783 & n13508 ;
  assign n13517 = n13510 | n13516 ;
  assign n10571 = n5838 & n10542 ;
  assign n10515 = x[122] & n10481 ;
  assign n11889 = x[123] & n11232 ;
  assign n13518 = n10515 | n11889 ;
  assign n13519 = x[124] & n10479 ;
  assign n13520 = n13518 | n13519 ;
  assign n13521 = n10571 | n13520 ;
  assign n31824 = ~n13521 ;
  assign n13522 = x[14] & n31824 ;
  assign n13523 = n27956 & n13521 ;
  assign n13524 = n13522 | n13523 ;
  assign n31825 = ~n13524 ;
  assign n13525 = n13517 & n31825 ;
  assign n31826 = ~n13517 ;
  assign n13526 = n31826 & n13524 ;
  assign n13527 = n13525 | n13526 ;
  assign n8743 = n4985 & n8706 ;
  assign n8689 = x[119] & n8645 ;
  assign n9863 = x[120] & n9278 ;
  assign n11959 = n8689 | n9863 ;
  assign n11960 = x[121] & n8643 ;
  assign n11961 = n11959 | n11960 ;
  assign n11962 = n8743 | n11961 ;
  assign n11963 = x[17] | n11962 ;
  assign n11964 = x[17] & n11962 ;
  assign n31827 = ~n11964 ;
  assign n11965 = n11963 & n31827 ;
  assign n12603 = n11972 & n12601 ;
  assign n12609 = n12605 & n12607 ;
  assign n12610 = n12603 | n12609 ;
  assign n31828 = ~n12610 ;
  assign n12611 = n11965 & n31828 ;
  assign n31829 = ~n11965 ;
  assign n12613 = n31829 & n12610 ;
  assign n12614 = n12611 | n12613 ;
  assign n11808 = n11797 & n11806 ;
  assign n11814 = n11810 & n11812 ;
  assign n11815 = n11808 | n11814 ;
  assign n7204 = n784 & n7162 ;
  assign n7120 = x[116] & n7100 ;
  assign n7721 = x[117] & n7647 ;
  assign n11816 = n7120 | n7721 ;
  assign n11817 = x[118] & n7098 ;
  assign n11818 = n11816 | n11817 ;
  assign n11819 = n7204 | n11818 ;
  assign n31830 = ~n11819 ;
  assign n11820 = x[20] & n31830 ;
  assign n11821 = n28114 & n11819 ;
  assign n11822 = n11820 | n11821 ;
  assign n11823 = n11815 | n11822 ;
  assign n11824 = n11815 & n11822 ;
  assign n31831 = ~n11824 ;
  assign n11825 = n11823 & n31831 ;
  assign n4443 = n452 & n4442 ;
  assign n378 = x[110] & n330 ;
  assign n406 = x[111] & n390 ;
  assign n9952 = n378 | n406 ;
  assign n9953 = x[112] & n322 ;
  assign n9954 = n9952 | n9953 ;
  assign n9955 = n4443 | n9954 ;
  assign n31832 = ~n9955 ;
  assign n9956 = x[26] & n31832 ;
  assign n9957 = n28342 & n9955 ;
  assign n9958 = n9956 | n9957 ;
  assign n10426 = n9965 & n10424 ;
  assign n10432 = n10426 | n10431 ;
  assign n10433 = n9958 | n10432 ;
  assign n10434 = n9958 & n10432 ;
  assign n31833 = ~n10434 ;
  assign n10435 = n10433 & n31833 ;
  assign n9744 = n9736 | n9743 ;
  assign n4667 = n3639 & n4632 ;
  assign n4529 = x[107] & n4514 ;
  assign n4591 = x[108] & n4572 ;
  assign n9745 = n4529 | n4591 ;
  assign n9746 = x[109] & n4504 ;
  assign n9747 = n9745 | n9746 ;
  assign n9748 = n4667 | n9747 ;
  assign n31834 = ~n9748 ;
  assign n9749 = x[29] & n31834 ;
  assign n9750 = n28483 & n9748 ;
  assign n9751 = n9749 | n9750 ;
  assign n9752 = n9744 | n9751 ;
  assign n9753 = n9744 & n9751 ;
  assign n31835 = ~n9753 ;
  assign n9754 = n9752 & n31835 ;
  assign n9187 = n8818 & n9185 ;
  assign n9193 = n9187 | n9192 ;
  assign n3229 = n779 & n3223 ;
  assign n682 = x[104] & n663 ;
  assign n731 = x[105] & n720 ;
  assign n9194 = n682 | n731 ;
  assign n9195 = x[106] & n652 ;
  assign n9196 = n9194 | n9195 ;
  assign n9197 = n3229 | n9196 ;
  assign n31836 = ~n9197 ;
  assign n9198 = x[32] & n31836 ;
  assign n9199 = n28658 & n9197 ;
  assign n9200 = n9198 | n9199 ;
  assign n9201 = n9193 | n9200 ;
  assign n9202 = n9193 & n9200 ;
  assign n31837 = ~n9202 ;
  assign n9203 = n9201 & n31837 ;
  assign n8052 = n7770 & n8050 ;
  assign n8062 = n8059 & n8061 ;
  assign n8064 = n8052 | n8062 ;
  assign n7537 = n7528 & n7535 ;
  assign n7538 = n7527 | n7537 ;
  assign n6975 = n6966 & n6973 ;
  assign n6976 = n6965 | n6975 ;
  assign n6043 = n6040 & n6042 ;
  assign n6055 = n6043 | n6054 ;
  assign n2022 = n1720 & n2007 ;
  assign n1915 = x[86] & n1866 ;
  assign n1983 = x[87] & n1931 ;
  assign n5936 = n1915 | n1983 ;
  assign n5937 = x[88] & n1862 ;
  assign n5938 = n5936 | n5937 ;
  assign n5939 = n2022 | n5938 ;
  assign n31838 = ~n5939 ;
  assign n5940 = x[50] & n31838 ;
  assign n5941 = n29865 & n5939 ;
  assign n5942 = n5940 | n5941 ;
  assign n1467 = n1003 & n1457 ;
  assign n1367 = x[80] & n1319 ;
  assign n1428 = x[81] & n1384 ;
  assign n3682 = n1367 | n1428 ;
  assign n3683 = x[82] & n1315 ;
  assign n3684 = n3682 | n3683 ;
  assign n3685 = n1467 | n3684 ;
  assign n3686 = x[56] | n3685 ;
  assign n3687 = x[56] & n3685 ;
  assign n31839 = ~n3687 ;
  assign n3688 = n3686 & n31839 ;
  assign n3315 = n3282 & n3303 ;
  assign n3317 = n3315 | n3316 ;
  assign n917 = x[74] & n900 ;
  assign n985 = x[75] & n949 ;
  assign n2744 = n917 | n985 ;
  assign n2745 = x[76] & n881 ;
  assign n2746 = n2744 | n2745 ;
  assign n2759 = n1006 & n2750 ;
  assign n2760 = n2746 | n2759 ;
  assign n31840 = ~n2760 ;
  assign n2761 = x[62] & n31840 ;
  assign n2762 = n30886 & n2760 ;
  assign n2763 = n2761 | n2762 ;
  assign n27692 = x[72] & n27215 ;
  assign n835 = x[73] & n805 ;
  assign n1758 = n27692 | n835 ;
  assign n1760 = x[8] | n1759 ;
  assign n1761 = x[8] & n1759 ;
  assign n31841 = ~n1761 ;
  assign n1762 = n1760 & n31841 ;
  assign n31842 = ~n1758 ;
  assign n1763 = n31842 & n1762 ;
  assign n31843 = ~n1762 ;
  assign n1764 = n1758 & n31843 ;
  assign n2741 = n1763 | n1764 ;
  assign n31844 = ~n2741 ;
  assign n2742 = n2740 & n31844 ;
  assign n31845 = ~n2740 ;
  assign n2764 = n31845 & n2741 ;
  assign n2765 = n2742 | n2764 ;
  assign n31846 = ~n2763 ;
  assign n2766 = n31846 & n2765 ;
  assign n31847 = ~n2765 ;
  assign n3268 = n2763 & n31847 ;
  assign n3269 = n2766 | n3268 ;
  assign n1747 = n1217 & n1741 ;
  assign n1114 = x[77] & n1079 ;
  assign n1165 = x[78] & n1144 ;
  assign n3270 = n1114 | n1165 ;
  assign n3271 = x[79] & n1075 ;
  assign n3272 = n3270 | n3271 ;
  assign n3273 = n1747 | n3272 ;
  assign n31848 = ~n3273 ;
  assign n3274 = x[59] & n31848 ;
  assign n3275 = n30638 & n3273 ;
  assign n3276 = n3274 | n3275 ;
  assign n3277 = n3269 | n3276 ;
  assign n3278 = n3269 & n3276 ;
  assign n31849 = ~n3278 ;
  assign n3318 = n3277 & n31849 ;
  assign n3319 = n3317 & n3318 ;
  assign n3689 = n3317 | n3318 ;
  assign n31850 = ~n3319 ;
  assign n3690 = n31850 & n3689 ;
  assign n3691 = n3688 & n3690 ;
  assign n3692 = n3688 | n3690 ;
  assign n31851 = ~n3691 ;
  assign n3693 = n31851 & n3692 ;
  assign n3780 = n3771 & n3778 ;
  assign n3781 = n3769 | n3780 ;
  assign n31852 = ~n3781 ;
  assign n3782 = n3693 & n31852 ;
  assign n31853 = ~n3693 ;
  assign n4755 = n31853 & n3781 ;
  assign n4756 = n3782 | n4755 ;
  assign n1697 = n1239 & n1690 ;
  assign n1597 = x[83] & n1551 ;
  assign n1660 = x[84] & n1616 ;
  assign n4757 = n1597 | n1660 ;
  assign n4758 = x[85] & n1547 ;
  assign n4759 = n4757 | n4758 ;
  assign n4760 = n1697 | n4759 ;
  assign n31854 = ~n4760 ;
  assign n4761 = x[53] & n31854 ;
  assign n4762 = n30125 & n4760 ;
  assign n4763 = n4761 | n4762 ;
  assign n31855 = ~n4763 ;
  assign n4764 = n4756 & n31855 ;
  assign n31856 = ~n4756 ;
  assign n4766 = n31856 & n4763 ;
  assign n4767 = n4764 | n4766 ;
  assign n4855 = n4846 & n4853 ;
  assign n4856 = n4845 | n4855 ;
  assign n31857 = ~n4856 ;
  assign n4857 = n4767 & n31857 ;
  assign n31858 = ~n4767 ;
  assign n5943 = n31858 & n4856 ;
  assign n5944 = n4857 | n5943 ;
  assign n31859 = ~n5942 ;
  assign n5945 = n31859 & n5944 ;
  assign n31860 = ~n5944 ;
  assign n6056 = n5942 & n31860 ;
  assign n6057 = n5945 | n6056 ;
  assign n6058 = n6055 | n6057 ;
  assign n6059 = n6055 & n6057 ;
  assign n31861 = ~n6059 ;
  assign n6344 = n6058 & n31861 ;
  assign n2330 = n2046 & n2321 ;
  assign n2202 = x[89] & n2179 ;
  assign n2291 = x[90] & n2244 ;
  assign n6345 = n2202 | n2291 ;
  assign n6346 = x[91] & n2175 ;
  assign n6347 = n6345 | n6346 ;
  assign n6348 = n2330 | n6347 ;
  assign n31862 = ~n6348 ;
  assign n6349 = x[47] & n31862 ;
  assign n6350 = n29621 & n6348 ;
  assign n6351 = n6349 | n6350 ;
  assign n31863 = ~n6351 ;
  assign n6352 = n6344 & n31863 ;
  assign n31864 = ~n6344 ;
  assign n6354 = n31864 & n6351 ;
  assign n6355 = n6352 | n6354 ;
  assign n6593 = n6591 & n6592 ;
  assign n6595 = n6584 | n6593 ;
  assign n31865 = ~n6595 ;
  assign n6596 = n6355 & n31865 ;
  assign n31866 = ~n6355 ;
  assign n6770 = n31866 & n6595 ;
  assign n6771 = n6596 | n6770 ;
  assign n2651 = n2410 & n2635 ;
  assign n2542 = x[92] & n2492 ;
  assign n2598 = x[93] & n2557 ;
  assign n6772 = n2542 | n2598 ;
  assign n6773 = x[94] & n2488 ;
  assign n6774 = n6772 | n6773 ;
  assign n6775 = n2651 | n6774 ;
  assign n31867 = ~n6775 ;
  assign n6776 = x[44] & n31867 ;
  assign n6777 = n29400 & n6775 ;
  assign n6778 = n6776 | n6777 ;
  assign n6779 = n6771 & n6778 ;
  assign n6977 = n6771 | n6778 ;
  assign n31868 = ~n6779 ;
  assign n7277 = n31868 & n6977 ;
  assign n31869 = ~n7277 ;
  assign n7278 = n6976 & n31869 ;
  assign n6978 = n6976 & n6977 ;
  assign n6979 = n6779 | n6978 ;
  assign n31870 = ~n6979 ;
  assign n7279 = n6977 & n31870 ;
  assign n7280 = n7278 | n7279 ;
  assign n3186 = n2438 & n3162 ;
  assign n3046 = x[95] & n3031 ;
  assign n3130 = x[96] & n3096 ;
  assign n7281 = n3046 | n3130 ;
  assign n7282 = x[97] & n3027 ;
  assign n7283 = n7281 | n7282 ;
  assign n7284 = n3186 | n7283 ;
  assign n31871 = ~n7284 ;
  assign n7285 = x[41] & n31871 ;
  assign n7286 = n29184 & n7284 ;
  assign n7287 = n7285 | n7286 ;
  assign n31872 = ~n7287 ;
  assign n7288 = n7280 & n31872 ;
  assign n31873 = ~n7280 ;
  assign n7539 = n31873 & n7287 ;
  assign n7540 = n7288 | n7539 ;
  assign n7541 = n7538 | n7540 ;
  assign n7542 = n7538 & n7540 ;
  assign n31874 = ~n7542 ;
  assign n7759 = n7541 & n31874 ;
  assign n3595 = n2466 & n3574 ;
  assign n3495 = x[98] & n3443 ;
  assign n3556 = x[99] & n3508 ;
  assign n7760 = n3495 | n3556 ;
  assign n7761 = x[100] & n3439 ;
  assign n7762 = n7760 | n7761 ;
  assign n7763 = n3595 | n7762 ;
  assign n31875 = ~n7763 ;
  assign n7764 = x[38] & n31875 ;
  assign n7765 = n28996 & n7763 ;
  assign n7766 = n7764 | n7765 ;
  assign n7767 = n7759 | n7766 ;
  assign n7768 = n7759 & n7766 ;
  assign n31876 = ~n7768 ;
  assign n8065 = n7767 & n31876 ;
  assign n31877 = ~n8064 ;
  assign n8066 = n31877 & n8065 ;
  assign n31878 = ~n8065 ;
  assign n8213 = n8064 & n31878 ;
  assign n8214 = n8066 | n8213 ;
  assign n4069 = n2626 & n4041 ;
  assign n3929 = x[101] & n3910 ;
  assign n4004 = x[102] & n3975 ;
  assign n8215 = n3929 | n4004 ;
  assign n8216 = x[103] & n3906 ;
  assign n8217 = n8215 | n8216 ;
  assign n8218 = n4069 | n8217 ;
  assign n31879 = ~n8218 ;
  assign n8219 = x[35] & n31879 ;
  assign n8220 = n28822 & n8218 ;
  assign n8221 = n8219 | n8220 ;
  assign n31880 = ~n8221 ;
  assign n8222 = n8214 & n31880 ;
  assign n31881 = ~n8214 ;
  assign n8224 = n31881 & n8221 ;
  assign n8225 = n8222 | n8224 ;
  assign n8556 = n8546 | n8555 ;
  assign n8557 = n8225 | n8556 ;
  assign n8558 = n8225 & n8556 ;
  assign n31882 = ~n8558 ;
  assign n9204 = n8557 & n31882 ;
  assign n31883 = ~n9204 ;
  assign n9205 = n9203 & n31883 ;
  assign n31884 = ~n9203 ;
  assign n9755 = n31884 & n9204 ;
  assign n9756 = n9205 | n9755 ;
  assign n31885 = ~n9756 ;
  assign n9758 = n9754 & n31885 ;
  assign n31886 = ~n9754 ;
  assign n10436 = n31886 & n9756 ;
  assign n10437 = n9758 | n10436 ;
  assign n31887 = ~n10437 ;
  assign n10438 = n10435 & n31887 ;
  assign n31888 = ~n10435 ;
  assign n11195 = n31888 & n10437 ;
  assign n11196 = n10438 | n11195 ;
  assign n5344 = n4474 & n5302 ;
  assign n5262 = x[113] & n5240 ;
  assign n6256 = x[114] & n6179 ;
  assign n10634 = n5262 | n6256 ;
  assign n10635 = x[115] & n5238 ;
  assign n10636 = n10634 | n10635 ;
  assign n10637 = n5344 | n10636 ;
  assign n31889 = ~n10637 ;
  assign n10638 = x[23] & n31889 ;
  assign n10639 = n28221 & n10637 ;
  assign n10640 = n10638 | n10639 ;
  assign n11186 = n10647 & n11184 ;
  assign n11191 = n11188 & n11189 ;
  assign n11192 = n11186 | n11191 ;
  assign n11193 = n10640 | n11192 ;
  assign n11194 = n10640 & n11192 ;
  assign n31890 = ~n11194 ;
  assign n11197 = n11193 & n31890 ;
  assign n11198 = n11196 & n11197 ;
  assign n11826 = n11196 | n11197 ;
  assign n31891 = ~n11198 ;
  assign n11827 = n31891 & n11826 ;
  assign n11828 = n11825 | n11827 ;
  assign n11829 = n11825 & n11827 ;
  assign n31892 = ~n11829 ;
  assign n12615 = n11828 & n31892 ;
  assign n12616 = n12614 & n12615 ;
  assign n13528 = n12614 | n12615 ;
  assign n13529 = n13527 & n13528 ;
  assign n31893 = ~n12616 ;
  assign n13530 = n31893 & n13529 ;
  assign n31894 = ~n13530 ;
  assign n14420 = n13527 & n31894 ;
  assign n14421 = n13528 & n31894 ;
  assign n14422 = n31893 & n14421 ;
  assign n14423 = n14420 | n14422 ;
  assign n31895 = ~n14423 ;
  assign n14424 = n14419 & n31895 ;
  assign n31896 = ~n14419 ;
  assign n15386 = n31896 & n14423 ;
  assign n15387 = n14424 | n15386 ;
  assign n15388 = n15385 | n15387 ;
  assign n15389 = n15385 & n15387 ;
  assign n31897 = ~n15389 ;
  assign n23139 = n15388 & n31897 ;
  assign n23140 = n23138 & n23139 ;
  assign n31898 = ~n15387 ;
  assign n27738 = n15385 & n31898 ;
  assign n31899 = ~n15385 ;
  assign n27739 = n31899 & n15387 ;
  assign n27740 = n23138 | n27739 ;
  assign n27741 = n27738 | n27740 ;
  assign n31900 = ~n23140 ;
  assign n201 = n31900 & n27741 ;
  assign n23141 = n15389 | n23140 ;
  assign n14425 = n14419 & n14423 ;
  assign n14426 = n14418 | n14425 ;
  assign n10576 = n642 & n10542 ;
  assign n10520 = x[123] & n10481 ;
  assign n11873 = x[124] & n11232 ;
  assign n11952 = n10520 | n11873 ;
  assign n11953 = x[125] & n10479 ;
  assign n11954 = n11952 | n11953 ;
  assign n11955 = n10576 | n11954 ;
  assign n31901 = ~n11955 ;
  assign n11956 = x[14] & n31901 ;
  assign n11957 = n27956 & n11955 ;
  assign n11958 = n11956 | n11957 ;
  assign n12612 = n11965 & n12610 ;
  assign n12617 = n12612 | n12616 ;
  assign n12618 = n11958 | n12617 ;
  assign n12619 = n11958 & n12617 ;
  assign n31902 = ~n12619 ;
  assign n12620 = n12618 & n31902 ;
  assign n7209 = n5047 & n7162 ;
  assign n7115 = x[117] & n7100 ;
  assign n7700 = x[118] & n7647 ;
  assign n10627 = n7115 | n7700 ;
  assign n10628 = x[119] & n7098 ;
  assign n10629 = n10627 | n10628 ;
  assign n10630 = n7209 | n10629 ;
  assign n10631 = x[20] | n10630 ;
  assign n10632 = x[20] & n10630 ;
  assign n31903 = ~n10632 ;
  assign n10633 = n10631 & n31903 ;
  assign n11199 = n11194 | n11198 ;
  assign n31904 = ~n11199 ;
  assign n11200 = n10633 & n31904 ;
  assign n31905 = ~n10633 ;
  assign n11202 = n31905 & n11199 ;
  assign n11203 = n11200 | n11202 ;
  assign n5305 = n4702 & n5302 ;
  assign n5267 = x[114] & n5240 ;
  assign n6257 = x[115] & n6179 ;
  assign n9945 = n5267 | n6257 ;
  assign n9946 = x[116] & n5238 ;
  assign n9947 = n9945 | n9946 ;
  assign n9948 = n5305 | n9947 ;
  assign n9949 = x[23] | n9948 ;
  assign n9950 = x[23] & n9948 ;
  assign n31906 = ~n9950 ;
  assign n9951 = n9949 & n31906 ;
  assign n10439 = n10435 & n10437 ;
  assign n10440 = n10434 | n10439 ;
  assign n31907 = ~n10440 ;
  assign n10441 = n9951 & n31907 ;
  assign n31908 = ~n9951 ;
  assign n10443 = n31908 & n10440 ;
  assign n10444 = n10441 | n10443 ;
  assign n4090 = n452 & n4087 ;
  assign n377 = x[111] & n330 ;
  assign n401 = x[112] & n390 ;
  assign n9301 = n377 | n401 ;
  assign n9302 = x[113] & n322 ;
  assign n9303 = n9301 | n9302 ;
  assign n9304 = n4090 | n9303 ;
  assign n31909 = ~n9304 ;
  assign n9305 = x[26] & n31909 ;
  assign n9306 = n28342 & n9304 ;
  assign n9307 = n9305 | n9306 ;
  assign n9757 = n9754 & n9756 ;
  assign n9759 = n9753 | n9757 ;
  assign n9760 = n9307 | n9759 ;
  assign n9761 = n9307 & n9759 ;
  assign n31910 = ~n9761 ;
  assign n9762 = n9760 & n31910 ;
  assign n3200 = n779 & n3199 ;
  assign n699 = x[105] & n663 ;
  assign n739 = x[106] & n720 ;
  assign n8206 = n699 | n739 ;
  assign n8207 = x[107] & n652 ;
  assign n8208 = n8206 | n8207 ;
  assign n8209 = n3200 | n8208 ;
  assign n31911 = ~n8209 ;
  assign n8210 = x[32] & n31911 ;
  assign n8211 = n28658 & n8209 ;
  assign n8212 = n8210 | n8211 ;
  assign n8223 = n8214 & n8221 ;
  assign n8559 = n8223 | n8558 ;
  assign n8560 = n8212 | n8559 ;
  assign n8561 = n8212 & n8559 ;
  assign n31912 = ~n8561 ;
  assign n8562 = n8560 & n31912 ;
  assign n4065 = n3001 & n4041 ;
  assign n3952 = x[102] & n3910 ;
  assign n4027 = x[103] & n3975 ;
  assign n8074 = n3952 | n4027 ;
  assign n8075 = x[104] & n3906 ;
  assign n8076 = n8074 | n8075 ;
  assign n8077 = n4065 | n8076 ;
  assign n8078 = x[35] | n8077 ;
  assign n8079 = x[35] & n8077 ;
  assign n31913 = ~n8079 ;
  assign n8080 = n8078 & n31913 ;
  assign n8067 = n8064 & n8065 ;
  assign n8068 = n7768 | n8067 ;
  assign n3605 = n2977 & n3574 ;
  assign n3475 = x[99] & n3443 ;
  assign n3554 = x[100] & n3508 ;
  assign n7547 = n3475 | n3554 ;
  assign n7548 = x[101] & n3439 ;
  assign n7549 = n7547 | n7548 ;
  assign n7550 = n3605 | n7549 ;
  assign n7551 = x[38] | n7550 ;
  assign n7552 = x[38] & n7550 ;
  assign n31914 = ~n7552 ;
  assign n7553 = n7551 & n31914 ;
  assign n7289 = n7280 & n7287 ;
  assign n7543 = n7289 | n7542 ;
  assign n3182 = n2841 & n3162 ;
  assign n3054 = x[96] & n3031 ;
  assign n3143 = x[97] & n3096 ;
  assign n6983 = n3054 | n3143 ;
  assign n6984 = x[98] & n3027 ;
  assign n6985 = n6983 | n6984 ;
  assign n6986 = n3182 | n6985 ;
  assign n6987 = x[41] | n6986 ;
  assign n6988 = x[41] & n6986 ;
  assign n31915 = ~n6988 ;
  assign n6989 = n6987 & n31915 ;
  assign n932 = x[75] & n900 ;
  assign n957 = x[76] & n949 ;
  assign n1769 = n932 | n957 ;
  assign n1770 = x[77] & n881 ;
  assign n1771 = n1769 | n1770 ;
  assign n1781 = n1006 & n1775 ;
  assign n1782 = n1771 | n1781 ;
  assign n31916 = ~n1782 ;
  assign n1783 = x[62] & n31916 ;
  assign n1784 = n30886 & n1782 ;
  assign n1785 = n1783 | n1784 ;
  assign n27679 = x[73] & n27215 ;
  assign n831 = x[74] & n805 ;
  assign n1253 = n27679 | n831 ;
  assign n1765 = n27845 & n1759 ;
  assign n1766 = n1764 | n1765 ;
  assign n1767 = n1253 | n1766 ;
  assign n1786 = n1253 & n1766 ;
  assign n31917 = ~n1786 ;
  assign n1787 = n1767 & n31917 ;
  assign n31918 = ~n1785 ;
  assign n1788 = n31918 & n1787 ;
  assign n31919 = ~n1787 ;
  assign n1789 = n1785 & n31919 ;
  assign n2702 = n1788 | n1789 ;
  assign n2743 = n2740 | n2741 ;
  assign n2767 = n2763 & n2765 ;
  assign n31920 = ~n2767 ;
  assign n2768 = n2743 & n31920 ;
  assign n31921 = ~n2702 ;
  assign n2769 = n31921 & n2768 ;
  assign n31922 = ~n2768 ;
  assign n2771 = n2702 & n31922 ;
  assign n2772 = n2769 | n2771 ;
  assign n1272 = n1217 & n1270 ;
  assign n1111 = x[78] & n1079 ;
  assign n1176 = x[79] & n1144 ;
  assign n2773 = n1111 | n1176 ;
  assign n2774 = x[80] & n1075 ;
  assign n2775 = n2773 | n2774 ;
  assign n2776 = n1272 | n2775 ;
  assign n31923 = ~n2776 ;
  assign n2777 = x[59] & n31923 ;
  assign n2778 = n30638 & n2776 ;
  assign n2779 = n2777 | n2778 ;
  assign n31924 = ~n2779 ;
  assign n2780 = n2772 & n31924 ;
  assign n31925 = ~n2772 ;
  assign n3266 = n31925 & n2779 ;
  assign n3267 = n2780 | n3266 ;
  assign n3320 = n3278 | n3319 ;
  assign n3321 = n3267 | n3320 ;
  assign n3322 = n3267 & n3320 ;
  assign n31926 = ~n3322 ;
  assign n3323 = n3321 & n31926 ;
  assign n1466 = n1057 & n1457 ;
  assign n1381 = x[81] & n1319 ;
  assign n1416 = x[82] & n1384 ;
  assign n3324 = n1381 | n1416 ;
  assign n3325 = x[83] & n1315 ;
  assign n3326 = n3324 | n3325 ;
  assign n3327 = n1466 | n3326 ;
  assign n31927 = ~n3327 ;
  assign n3328 = x[56] & n31927 ;
  assign n3329 = n30379 & n3327 ;
  assign n3330 = n3328 | n3329 ;
  assign n31928 = ~n3330 ;
  assign n3331 = n3323 & n31928 ;
  assign n31929 = ~n3323 ;
  assign n3680 = n31929 & n3330 ;
  assign n3681 = n3331 | n3680 ;
  assign n3783 = n3693 & n3781 ;
  assign n3784 = n3691 | n3783 ;
  assign n3785 = n3681 | n3784 ;
  assign n3786 = n3681 & n3784 ;
  assign n31930 = ~n3786 ;
  assign n3787 = n3785 & n31930 ;
  assign n1693 = n1213 & n1690 ;
  assign n1595 = x[84] & n1551 ;
  assign n1618 = x[85] & n1616 ;
  assign n3788 = n1595 | n1618 ;
  assign n3789 = x[86] & n1547 ;
  assign n3790 = n3788 | n3789 ;
  assign n3791 = n1693 | n3790 ;
  assign n31931 = ~n3791 ;
  assign n3792 = x[53] & n31931 ;
  assign n3793 = n30125 & n3791 ;
  assign n3794 = n3792 | n3793 ;
  assign n31932 = ~n3794 ;
  assign n3795 = n3787 & n31932 ;
  assign n31933 = ~n3787 ;
  assign n4753 = n31933 & n3794 ;
  assign n4754 = n3795 | n4753 ;
  assign n4765 = n4756 & n4763 ;
  assign n4858 = n4767 & n4856 ;
  assign n4859 = n4765 | n4858 ;
  assign n4860 = n4754 | n4859 ;
  assign n4861 = n4754 & n4859 ;
  assign n31934 = ~n4861 ;
  assign n4862 = n4860 & n31934 ;
  assign n2014 = n1453 & n2007 ;
  assign n1926 = x[87] & n1866 ;
  assign n1963 = x[88] & n1931 ;
  assign n4863 = n1926 | n1963 ;
  assign n4864 = x[89] & n1862 ;
  assign n4865 = n4863 | n4864 ;
  assign n4866 = n2014 | n4865 ;
  assign n31935 = ~n4866 ;
  assign n4867 = x[50] & n31935 ;
  assign n4868 = n29865 & n4866 ;
  assign n4869 = n4867 | n4868 ;
  assign n31936 = ~n4869 ;
  assign n4870 = n4862 & n31936 ;
  assign n31937 = ~n4862 ;
  assign n5934 = n31937 & n4869 ;
  assign n5935 = n4870 | n5934 ;
  assign n5946 = n5942 & n5944 ;
  assign n6060 = n5946 | n6059 ;
  assign n6061 = n5935 | n6060 ;
  assign n6062 = n5935 & n6060 ;
  assign n31938 = ~n6062 ;
  assign n6063 = n6061 & n31938 ;
  assign n2337 = n1841 & n2321 ;
  assign n2190 = x[90] & n2179 ;
  assign n2289 = x[91] & n2244 ;
  assign n6064 = n2190 | n2289 ;
  assign n6065 = x[92] & n2175 ;
  assign n6066 = n6064 | n6065 ;
  assign n6067 = n2337 | n6066 ;
  assign n31939 = ~n6067 ;
  assign n6068 = x[47] & n31939 ;
  assign n6069 = n29621 & n6067 ;
  assign n6070 = n6068 | n6069 ;
  assign n31940 = ~n6070 ;
  assign n6071 = n6063 & n31940 ;
  assign n31941 = ~n6063 ;
  assign n6342 = n31941 & n6070 ;
  assign n6343 = n6071 | n6342 ;
  assign n6353 = n6344 & n6351 ;
  assign n6597 = n6355 & n6595 ;
  assign n6598 = n6353 | n6597 ;
  assign n31942 = ~n6598 ;
  assign n6599 = n6343 & n31942 ;
  assign n31943 = ~n6343 ;
  assign n6601 = n31943 & n6598 ;
  assign n6602 = n6599 | n6601 ;
  assign n2650 = n2152 & n2635 ;
  assign n2528 = x[93] & n2492 ;
  assign n2590 = x[94] & n2557 ;
  assign n6603 = n2528 | n2590 ;
  assign n6604 = x[95] & n2488 ;
  assign n6605 = n6603 | n6604 ;
  assign n6606 = n2650 | n6605 ;
  assign n31944 = ~n6606 ;
  assign n6607 = x[44] & n31944 ;
  assign n6608 = n29400 & n6606 ;
  assign n6609 = n6607 | n6608 ;
  assign n31945 = ~n6609 ;
  assign n6610 = n6602 & n31945 ;
  assign n31946 = ~n6602 ;
  assign n6980 = n31946 & n6609 ;
  assign n6981 = n6610 | n6980 ;
  assign n6982 = n6979 & n6981 ;
  assign n6990 = n6979 | n6981 ;
  assign n31947 = ~n6982 ;
  assign n6991 = n31947 & n6990 ;
  assign n6992 = n6989 & n6991 ;
  assign n7544 = n6989 | n6991 ;
  assign n31948 = ~n6992 ;
  assign n7545 = n31948 & n7544 ;
  assign n31949 = ~n7545 ;
  assign n7554 = n7543 & n31949 ;
  assign n31950 = ~n7543 ;
  assign n7555 = n31950 & n7545 ;
  assign n7556 = n7554 | n7555 ;
  assign n7557 = n7553 & n7556 ;
  assign n8069 = n7553 | n7555 ;
  assign n8070 = n7554 | n8069 ;
  assign n31951 = ~n7557 ;
  assign n8071 = n31951 & n8070 ;
  assign n8072 = n8068 | n8071 ;
  assign n8073 = n8068 & n8071 ;
  assign n31952 = ~n8073 ;
  assign n8081 = n8072 & n31952 ;
  assign n31953 = ~n8081 ;
  assign n8082 = n8080 & n31953 ;
  assign n31954 = ~n8080 ;
  assign n8563 = n31954 & n8081 ;
  assign n8564 = n8082 | n8563 ;
  assign n31955 = ~n8564 ;
  assign n8565 = n8562 & n31955 ;
  assign n31956 = ~n8562 ;
  assign n9219 = n31956 & n8564 ;
  assign n9220 = n8565 | n9219 ;
  assign n9206 = n9203 & n9204 ;
  assign n9207 = n9202 | n9206 ;
  assign n4507 = x[110] & n4504 ;
  assign n9208 = x[108] & n4514 ;
  assign n9209 = x[109] & n4572 ;
  assign n9210 = n9208 | n9209 ;
  assign n9211 = n4507 | n9210 ;
  assign n9212 = n3615 & n4632 ;
  assign n9213 = n9211 | n9212 ;
  assign n9214 = n28483 & n9213 ;
  assign n31957 = ~n9213 ;
  assign n9215 = x[29] & n31957 ;
  assign n9216 = n9214 | n9215 ;
  assign n31958 = ~n9216 ;
  assign n9217 = n9207 & n31958 ;
  assign n31959 = ~n9207 ;
  assign n9221 = n31959 & n9216 ;
  assign n9222 = n9217 | n9221 ;
  assign n31960 = ~n9222 ;
  assign n9223 = n9220 & n31960 ;
  assign n31961 = ~n9220 ;
  assign n9763 = n31961 & n9222 ;
  assign n9764 = n9223 | n9763 ;
  assign n9765 = n9762 | n9764 ;
  assign n9766 = n9762 & n9764 ;
  assign n31962 = ~n9766 ;
  assign n10445 = n9765 & n31962 ;
  assign n10446 = n10444 & n10445 ;
  assign n11204 = n10444 | n10445 ;
  assign n11205 = n11203 & n11204 ;
  assign n31963 = ~n10446 ;
  assign n11206 = n31963 & n11205 ;
  assign n31964 = ~n11206 ;
  assign n11207 = n11203 & n31964 ;
  assign n11842 = n11204 & n31964 ;
  assign n11843 = n31963 & n11842 ;
  assign n11844 = n11207 | n11843 ;
  assign n11830 = n11824 | n11829 ;
  assign n9822 = x[122] & n8643 ;
  assign n11831 = x[120] & n8645 ;
  assign n11832 = x[121] & n9278 ;
  assign n11833 = n11831 | n11832 ;
  assign n11834 = n9822 | n11833 ;
  assign n11835 = n5022 & n8706 ;
  assign n11836 = n11834 | n11835 ;
  assign n11837 = n28039 & n11836 ;
  assign n31965 = ~n11836 ;
  assign n11838 = x[17] & n31965 ;
  assign n11839 = n11837 | n11838 ;
  assign n31966 = ~n11839 ;
  assign n11840 = n11830 & n31966 ;
  assign n31967 = ~n11830 ;
  assign n11845 = n31967 & n11839 ;
  assign n11846 = n11840 | n11845 ;
  assign n11847 = n11844 | n11846 ;
  assign n11848 = n11844 & n11846 ;
  assign n31968 = ~n11848 ;
  assign n12621 = n11847 & n31968 ;
  assign n31969 = ~n12621 ;
  assign n12622 = n12620 & n31969 ;
  assign n31970 = ~n12620 ;
  assign n13543 = n31970 & n12621 ;
  assign n13544 = n12622 | n13543 ;
  assign n13531 = n13517 & n13524 ;
  assign n13532 = n13530 | n13531 ;
  assign n12726 = n6186 & n12695 ;
  assign n13534 = x[126] & n12633 ;
  assign n13535 = x[127] & n13533 ;
  assign n13536 = n13534 | n13535 ;
  assign n13537 = n12726 | n13536 ;
  assign n31971 = ~n13537 ;
  assign n13538 = x[11] & n31971 ;
  assign n13539 = n27892 & n13537 ;
  assign n13540 = n13538 | n13539 ;
  assign n31972 = ~n13540 ;
  assign n13541 = n13532 & n31972 ;
  assign n31973 = ~n13532 ;
  assign n13545 = n31973 & n13540 ;
  assign n13546 = n13541 | n13545 ;
  assign n13547 = n13544 & n13546 ;
  assign n14427 = n13544 | n13545 ;
  assign n14428 = n13541 | n14427 ;
  assign n31974 = ~n13547 ;
  assign n14429 = n31974 & n14428 ;
  assign n14430 = n14426 | n14429 ;
  assign n14431 = n14426 & n14429 ;
  assign n31975 = ~n14431 ;
  assign n23142 = n14430 & n31975 ;
  assign n23143 = n23141 & n23142 ;
  assign n31976 = ~n14429 ;
  assign n27743 = n14426 & n31976 ;
  assign n31977 = ~n14426 ;
  assign n27744 = n31977 & n14429 ;
  assign n27745 = n23141 | n27744 ;
  assign n27746 = n27743 | n27745 ;
  assign n31978 = ~n23143 ;
  assign n202 = n31978 & n27746 ;
  assign n23144 = n14431 | n23143 ;
  assign n13542 = n13532 & n13540 ;
  assign n13548 = n13542 | n13547 ;
  assign n12623 = n12620 & n12621 ;
  assign n12624 = n12619 | n12623 ;
  assign n12676 = x[127] & n12633 ;
  assign n12734 = n5360 & n12695 ;
  assign n12759 = n12676 | n12734 ;
  assign n31979 = ~n12759 ;
  assign n12760 = x[11] & n31979 ;
  assign n12761 = n27892 & n12759 ;
  assign n12762 = n12760 | n12761 ;
  assign n12763 = n12624 | n12762 ;
  assign n12764 = n12624 & n12762 ;
  assign n31980 = ~n12764 ;
  assign n12765 = n12763 & n31980 ;
  assign n11841 = n11830 & n11839 ;
  assign n11849 = n11841 | n11848 ;
  assign n11850 = x[126] & n10479 ;
  assign n11853 = x[124] & n10481 ;
  assign n11854 = x[125] & n11232 ;
  assign n11855 = n11853 | n11854 ;
  assign n11856 = n11850 | n11855 ;
  assign n11857 = n5388 & n10542 ;
  assign n11858 = n11856 | n11857 ;
  assign n11859 = n27956 & n11858 ;
  assign n31981 = ~n11858 ;
  assign n11860 = x[14] & n31981 ;
  assign n11861 = n11859 | n11860 ;
  assign n31982 = ~n11861 ;
  assign n11862 = n11849 & n31982 ;
  assign n31983 = ~n11849 ;
  assign n11864 = n31983 & n11861 ;
  assign n11865 = n11862 | n11864 ;
  assign n8747 = n5417 & n8706 ;
  assign n8696 = x[121] & n8645 ;
  assign n9861 = x[122] & n9278 ;
  assign n10620 = n8696 | n9861 ;
  assign n10621 = x[123] & n8643 ;
  assign n10622 = n10620 | n10621 ;
  assign n10623 = n8747 | n10622 ;
  assign n31984 = ~n10623 ;
  assign n10624 = x[17] & n31984 ;
  assign n10625 = n28039 & n10623 ;
  assign n10626 = n10624 | n10625 ;
  assign n11201 = n10633 & n11199 ;
  assign n11208 = n11201 | n11206 ;
  assign n31985 = ~n11208 ;
  assign n11209 = n10626 & n31985 ;
  assign n31986 = ~n10626 ;
  assign n11211 = n31986 & n11208 ;
  assign n11212 = n11209 | n11211 ;
  assign n7190 = n4678 & n7162 ;
  assign n7146 = x[118] & n7100 ;
  assign n7709 = x[119] & n7647 ;
  assign n9938 = n7146 | n7709 ;
  assign n9939 = x[120] & n7098 ;
  assign n9940 = n9938 | n9939 ;
  assign n9941 = n7190 | n9940 ;
  assign n31987 = ~n9941 ;
  assign n9942 = x[20] & n31987 ;
  assign n9943 = n28114 & n9941 ;
  assign n9944 = n9942 | n9943 ;
  assign n10442 = n9951 & n10440 ;
  assign n10447 = n10442 | n10446 ;
  assign n10448 = n9944 | n10447 ;
  assign n10449 = n9944 & n10447 ;
  assign n31988 = ~n10449 ;
  assign n10450 = n10448 & n31988 ;
  assign n9218 = n9207 & n9216 ;
  assign n9224 = n9220 & n9222 ;
  assign n9225 = n9218 | n9224 ;
  assign n324 = x[114] & n322 ;
  assign n9226 = x[112] & n330 ;
  assign n9227 = x[113] & n390 ;
  assign n9228 = n9226 | n9227 ;
  assign n9229 = n324 | n9228 ;
  assign n9230 = n452 & n4276 ;
  assign n9231 = n9229 | n9230 ;
  assign n9232 = n28342 & n9231 ;
  assign n31989 = ~n9231 ;
  assign n9233 = x[26] & n31989 ;
  assign n9234 = n9232 | n9233 ;
  assign n31990 = ~n9234 ;
  assign n9235 = n9225 & n31990 ;
  assign n31991 = ~n9225 ;
  assign n9237 = n31991 & n9234 ;
  assign n9238 = n9235 | n9237 ;
  assign n4651 = n4246 & n4632 ;
  assign n4535 = x[109] & n4514 ;
  assign n4593 = x[110] & n4572 ;
  assign n8199 = n4535 | n4593 ;
  assign n8200 = x[111] & n4504 ;
  assign n8201 = n8199 | n8200 ;
  assign n8202 = n4651 | n8201 ;
  assign n31992 = ~n8202 ;
  assign n8203 = x[29] & n31992 ;
  assign n8204 = n28483 & n8202 ;
  assign n8205 = n8203 | n8204 ;
  assign n8566 = n8562 & n8564 ;
  assign n8567 = n8561 | n8566 ;
  assign n31993 = ~n8567 ;
  assign n8568 = n8205 & n31993 ;
  assign n31994 = ~n8205 ;
  assign n8570 = n31994 & n8567 ;
  assign n8571 = n8568 | n8570 ;
  assign n8083 = n8080 & n8081 ;
  assign n8084 = n8073 | n8083 ;
  assign n656 = x[108] & n652 ;
  assign n8085 = x[106] & n663 ;
  assign n8086 = x[107] & n720 ;
  assign n8087 = n8085 | n8086 ;
  assign n8088 = n656 | n8087 ;
  assign n8089 = n779 & n3876 ;
  assign n8090 = n8088 | n8089 ;
  assign n8091 = n28658 & n8090 ;
  assign n31995 = ~n8090 ;
  assign n8092 = x[32] & n31995 ;
  assign n8093 = n8091 | n8092 ;
  assign n8094 = n8084 | n8093 ;
  assign n8095 = n8084 & n8093 ;
  assign n31996 = ~n8095 ;
  assign n8096 = n8094 & n31996 ;
  assign n4078 = n3409 & n4041 ;
  assign n3950 = x[103] & n3910 ;
  assign n4026 = x[104] & n3975 ;
  assign n7563 = n3950 | n4026 ;
  assign n7564 = x[105] & n3906 ;
  assign n7565 = n7563 | n7564 ;
  assign n7566 = n4078 | n7565 ;
  assign n31997 = ~n7566 ;
  assign n7567 = x[35] & n31997 ;
  assign n7568 = n28822 & n7566 ;
  assign n7569 = n7567 | n7568 ;
  assign n7546 = n7543 & n7545 ;
  assign n7558 = n7546 | n7557 ;
  assign n3189 = n2313 & n3162 ;
  assign n3071 = x[97] & n3031 ;
  assign n3127 = x[98] & n3096 ;
  assign n6615 = n3071 | n3127 ;
  assign n6616 = x[99] & n3027 ;
  assign n6617 = n6615 | n6616 ;
  assign n6618 = n3189 | n6617 ;
  assign n31998 = ~n6618 ;
  assign n6619 = x[41] & n31998 ;
  assign n6620 = n29184 & n6618 ;
  assign n6621 = n6619 | n6620 ;
  assign n4871 = n4862 & n4869 ;
  assign n4872 = n4861 | n4871 ;
  assign n2011 = n1482 & n2007 ;
  assign n1898 = x[88] & n1866 ;
  assign n1964 = x[89] & n1931 ;
  assign n3803 = n1898 | n1964 ;
  assign n3804 = x[90] & n1862 ;
  assign n3805 = n3803 | n3804 ;
  assign n3806 = n2011 | n3805 ;
  assign n31999 = ~n3806 ;
  assign n3807 = x[50] & n31999 ;
  assign n3808 = n29865 & n3806 ;
  assign n3809 = n3807 | n3808 ;
  assign n3796 = n3787 & n3794 ;
  assign n3797 = n3786 | n3796 ;
  assign n1703 = n1522 & n1690 ;
  assign n1606 = x[85] & n1551 ;
  assign n1653 = x[86] & n1616 ;
  assign n3338 = n1606 | n1653 ;
  assign n3339 = x[87] & n1547 ;
  assign n3340 = n3338 | n3339 ;
  assign n3341 = n1703 | n3340 ;
  assign n3342 = x[53] | n3341 ;
  assign n3343 = x[53] & n3341 ;
  assign n32000 = ~n3343 ;
  assign n3344 = n3342 & n32000 ;
  assign n3332 = n3323 & n3330 ;
  assign n3333 = n3322 | n3332 ;
  assign n32001 = ~n1253 ;
  assign n1768 = n32001 & n1766 ;
  assign n1790 = n1768 | n1789 ;
  assign n27691 = x[74] & n27215 ;
  assign n833 = x[75] & n805 ;
  assign n1755 = n27691 | n833 ;
  assign n1756 = n1253 | n1755 ;
  assign n1791 = n1253 & n1755 ;
  assign n32002 = ~n1791 ;
  assign n1792 = n1756 & n32002 ;
  assign n32003 = ~n1790 ;
  assign n1793 = n32003 & n1792 ;
  assign n32004 = ~n1792 ;
  assign n1794 = n1790 & n32004 ;
  assign n2077 = n1793 | n1794 ;
  assign n929 = x[76] & n900 ;
  assign n981 = x[77] & n949 ;
  assign n2078 = n929 | n981 ;
  assign n2079 = x[78] & n881 ;
  assign n2080 = n2078 | n2079 ;
  assign n2091 = n1006 & n2084 ;
  assign n2092 = n2080 | n2091 ;
  assign n32005 = ~n2092 ;
  assign n2093 = x[62] & n32005 ;
  assign n2094 = n30886 & n2092 ;
  assign n2095 = n2093 | n2094 ;
  assign n32006 = ~n2095 ;
  assign n2096 = n2077 & n32006 ;
  assign n32007 = ~n2077 ;
  assign n2097 = n32007 & n2095 ;
  assign n2098 = n2096 | n2097 ;
  assign n1219 = n1029 & n1217 ;
  assign n1089 = x[79] & n1079 ;
  assign n1192 = x[80] & n1144 ;
  assign n2099 = n1089 | n1192 ;
  assign n2100 = x[81] & n1075 ;
  assign n2101 = n2099 | n2100 ;
  assign n2102 = n1219 | n2101 ;
  assign n32008 = ~n2102 ;
  assign n2103 = x[59] & n32008 ;
  assign n2104 = n30638 & n2102 ;
  assign n2105 = n2103 | n2104 ;
  assign n32009 = ~n2105 ;
  assign n2106 = n2098 & n32009 ;
  assign n32010 = ~n2098 ;
  assign n2107 = n32010 & n2105 ;
  assign n2701 = n2106 | n2107 ;
  assign n2770 = n2702 | n2768 ;
  assign n2781 = n2772 & n2779 ;
  assign n32011 = ~n2781 ;
  assign n2782 = n2770 & n32011 ;
  assign n2783 = n2701 & n2782 ;
  assign n2784 = n2701 | n2782 ;
  assign n32012 = ~n2783 ;
  assign n2785 = n32012 & n2784 ;
  assign n1465 = n1293 & n1457 ;
  assign n1350 = x[82] & n1319 ;
  assign n1414 = x[83] & n1384 ;
  assign n2786 = n1350 | n1414 ;
  assign n2787 = x[84] & n1315 ;
  assign n2788 = n2786 | n2787 ;
  assign n2789 = n1465 | n2788 ;
  assign n32013 = ~n2789 ;
  assign n2790 = x[56] & n32013 ;
  assign n2791 = n30379 & n2789 ;
  assign n2792 = n2790 | n2791 ;
  assign n32014 = ~n2792 ;
  assign n2793 = n2785 & n32014 ;
  assign n32015 = ~n2785 ;
  assign n3334 = n32015 & n2792 ;
  assign n3335 = n2793 | n3334 ;
  assign n32016 = ~n3333 ;
  assign n3336 = n32016 & n3335 ;
  assign n32017 = ~n3335 ;
  assign n3345 = n3333 & n32017 ;
  assign n3346 = n3336 | n3345 ;
  assign n3347 = n3344 & n3346 ;
  assign n3798 = n3336 | n3344 ;
  assign n3799 = n3345 | n3798 ;
  assign n32018 = ~n3347 ;
  assign n3800 = n32018 & n3799 ;
  assign n3801 = n3797 | n3800 ;
  assign n3802 = n3797 & n3800 ;
  assign n32019 = ~n3802 ;
  assign n3810 = n3801 & n32019 ;
  assign n3811 = n3809 & n3810 ;
  assign n4873 = n3809 | n3810 ;
  assign n32020 = ~n3811 ;
  assign n4874 = n32020 & n4873 ;
  assign n32021 = ~n4872 ;
  assign n4875 = n32021 & n4874 ;
  assign n32022 = ~n4874 ;
  assign n4877 = n4872 & n32022 ;
  assign n4878 = n4875 | n4877 ;
  assign n2341 = n1685 & n2321 ;
  assign n2224 = x[91] & n2179 ;
  assign n2277 = x[92] & n2244 ;
  assign n4879 = n2224 | n2277 ;
  assign n4880 = x[93] & n2175 ;
  assign n4881 = n4879 | n4880 ;
  assign n4882 = n2341 | n4881 ;
  assign n32023 = ~n4882 ;
  assign n4883 = x[47] & n32023 ;
  assign n4884 = n29621 & n4882 ;
  assign n4885 = n4883 | n4884 ;
  assign n32024 = ~n4885 ;
  assign n4886 = n4878 & n32024 ;
  assign n32025 = ~n4878 ;
  assign n5932 = n32025 & n4885 ;
  assign n5933 = n4886 | n5932 ;
  assign n6072 = n6063 & n6070 ;
  assign n6073 = n6062 | n6072 ;
  assign n6074 = n5933 | n6073 ;
  assign n6075 = n5933 & n6073 ;
  assign n32026 = ~n6075 ;
  assign n6076 = n6074 & n32026 ;
  assign n2648 = n2000 & n2635 ;
  assign n2517 = x[94] & n2492 ;
  assign n2606 = x[95] & n2557 ;
  assign n6077 = n2517 | n2606 ;
  assign n6078 = x[96] & n2488 ;
  assign n6079 = n6077 | n6078 ;
  assign n6080 = n2648 | n6079 ;
  assign n32027 = ~n6080 ;
  assign n6081 = x[44] & n32027 ;
  assign n6082 = n29400 & n6080 ;
  assign n6083 = n6081 | n6082 ;
  assign n32028 = ~n6083 ;
  assign n6084 = n6076 & n32028 ;
  assign n32029 = ~n6076 ;
  assign n6340 = n32029 & n6083 ;
  assign n6341 = n6084 | n6340 ;
  assign n6600 = n6343 & n6598 ;
  assign n6611 = n6602 & n6609 ;
  assign n6612 = n6600 | n6611 ;
  assign n32030 = ~n6612 ;
  assign n6613 = n6341 & n32030 ;
  assign n32031 = ~n6341 ;
  assign n6622 = n32031 & n6612 ;
  assign n6623 = n6613 | n6622 ;
  assign n32032 = ~n6621 ;
  assign n6624 = n32032 & n6623 ;
  assign n32033 = ~n6623 ;
  assign n6768 = n6621 & n32033 ;
  assign n6769 = n6624 | n6768 ;
  assign n6993 = n6982 | n6992 ;
  assign n6994 = n6769 | n6993 ;
  assign n6995 = n6769 & n6993 ;
  assign n32034 = ~n6995 ;
  assign n6996 = n6994 & n32034 ;
  assign n3601 = n2867 & n3574 ;
  assign n3482 = x[100] & n3443 ;
  assign n3546 = x[101] & n3508 ;
  assign n6997 = n3482 | n3546 ;
  assign n6998 = x[102] & n3439 ;
  assign n6999 = n6997 | n6998 ;
  assign n7000 = n3601 | n6999 ;
  assign n32035 = ~n7000 ;
  assign n7001 = x[38] & n32035 ;
  assign n7002 = n28996 & n7000 ;
  assign n7003 = n7001 | n7002 ;
  assign n32036 = ~n7003 ;
  assign n7004 = n6996 & n32036 ;
  assign n32037 = ~n6996 ;
  assign n7559 = n32037 & n7003 ;
  assign n7560 = n7004 | n7559 ;
  assign n32038 = ~n7558 ;
  assign n7561 = n32038 & n7560 ;
  assign n32039 = ~n7560 ;
  assign n7570 = n7558 & n32039 ;
  assign n7571 = n7561 | n7570 ;
  assign n32040 = ~n7569 ;
  assign n7572 = n32040 & n7571 ;
  assign n32041 = ~n7571 ;
  assign n8097 = n7569 & n32041 ;
  assign n8098 = n7572 | n8097 ;
  assign n32042 = ~n8098 ;
  assign n8099 = n8096 & n32042 ;
  assign n32043 = ~n8096 ;
  assign n8572 = n32043 & n8098 ;
  assign n8573 = n8099 | n8572 ;
  assign n8575 = n8571 & n8573 ;
  assign n8574 = n8571 | n8573 ;
  assign n9239 = n8574 & n9238 ;
  assign n32044 = ~n8575 ;
  assign n9240 = n32044 & n9239 ;
  assign n32045 = ~n9240 ;
  assign n9779 = n9238 & n32045 ;
  assign n9780 = n8574 & n32045 ;
  assign n9781 = n32044 & n9780 ;
  assign n9782 = n9779 | n9781 ;
  assign n9767 = n9761 | n9766 ;
  assign n6221 = x[117] & n5238 ;
  assign n9768 = x[115] & n5240 ;
  assign n9769 = x[116] & n6179 ;
  assign n9770 = n9768 | n9769 ;
  assign n9771 = n6221 | n9770 ;
  assign n9772 = n797 & n5302 ;
  assign n9773 = n9771 | n9772 ;
  assign n9774 = n28221 & n9773 ;
  assign n32046 = ~n9773 ;
  assign n9775 = x[23] & n32046 ;
  assign n9776 = n9774 | n9775 ;
  assign n32047 = ~n9776 ;
  assign n9777 = n9767 & n32047 ;
  assign n32048 = ~n9767 ;
  assign n9783 = n32048 & n9776 ;
  assign n9784 = n9777 | n9783 ;
  assign n9785 = n9782 | n9784 ;
  assign n9786 = n9782 & n9784 ;
  assign n32049 = ~n9786 ;
  assign n10451 = n9785 & n32049 ;
  assign n32050 = ~n10451 ;
  assign n10452 = n10450 & n32050 ;
  assign n32051 = ~n10450 ;
  assign n11213 = n32051 & n10451 ;
  assign n11214 = n10452 | n11213 ;
  assign n11216 = n11212 & n11214 ;
  assign n11215 = n11212 | n11214 ;
  assign n11867 = n11215 & n11865 ;
  assign n32052 = ~n11216 ;
  assign n11868 = n32052 & n11867 ;
  assign n32053 = ~n11868 ;
  assign n12766 = n11865 & n32053 ;
  assign n11866 = n32052 & n11865 ;
  assign n32054 = ~n11866 ;
  assign n12767 = n11215 & n32054 ;
  assign n12768 = n32052 & n12767 ;
  assign n12769 = n12766 | n12768 ;
  assign n32055 = ~n12769 ;
  assign n12770 = n12765 & n32055 ;
  assign n32056 = ~n12765 ;
  assign n13549 = n32056 & n12769 ;
  assign n13550 = n12770 | n13549 ;
  assign n13551 = n13548 | n13550 ;
  assign n13552 = n13548 & n13550 ;
  assign n32057 = ~n13552 ;
  assign n23145 = n13551 & n32057 ;
  assign n23146 = n23144 & n23145 ;
  assign n32058 = ~n13550 ;
  assign n27748 = n13548 & n32058 ;
  assign n32059 = ~n13548 ;
  assign n27749 = n32059 & n13550 ;
  assign n27750 = n23144 | n27749 ;
  assign n27751 = n27748 | n27750 ;
  assign n32060 = ~n23146 ;
  assign n203 = n32060 & n27751 ;
  assign n23147 = n13552 | n23146 ;
  assign n12771 = n12765 & n12769 ;
  assign n12772 = n12764 | n12771 ;
  assign n11863 = n11849 & n11861 ;
  assign n11869 = n11863 | n11868 ;
  assign n10580 = n5629 & n10542 ;
  assign n10523 = x[125] & n10481 ;
  assign n11892 = x[126] & n11232 ;
  assign n11929 = n10523 | n11892 ;
  assign n11930 = x[127] & n10479 ;
  assign n11931 = n11929 | n11930 ;
  assign n11932 = n10580 | n11931 ;
  assign n32061 = ~n11932 ;
  assign n11933 = x[14] & n32061 ;
  assign n11934 = n27956 & n11932 ;
  assign n11935 = n11933 | n11934 ;
  assign n11936 = n11869 | n11935 ;
  assign n11937 = n11869 & n11935 ;
  assign n32062 = ~n11937 ;
  assign n11938 = n11936 & n32062 ;
  assign n11210 = n10626 & n11208 ;
  assign n11217 = n11210 | n11216 ;
  assign n8718 = n5838 & n8706 ;
  assign n8674 = x[122] & n8645 ;
  assign n9864 = x[123] & n9278 ;
  assign n11218 = n8674 | n9864 ;
  assign n11219 = x[124] & n8643 ;
  assign n11220 = n11218 | n11219 ;
  assign n11221 = n8718 | n11220 ;
  assign n32063 = ~n11221 ;
  assign n11222 = x[17] & n32063 ;
  assign n11223 = n28039 & n11221 ;
  assign n11224 = n11222 | n11223 ;
  assign n11225 = n11217 | n11224 ;
  assign n11226 = n11217 & n11224 ;
  assign n32064 = ~n11226 ;
  assign n11227 = n11225 & n32064 ;
  assign n7206 = n4985 & n7162 ;
  assign n7124 = x[119] & n7100 ;
  assign n7684 = x[120] & n7647 ;
  assign n9931 = n7124 | n7684 ;
  assign n9932 = x[121] & n7098 ;
  assign n9933 = n9931 | n9932 ;
  assign n9934 = n7206 | n9933 ;
  assign n32065 = ~n9934 ;
  assign n9935 = x[20] & n32065 ;
  assign n9936 = n28114 & n9934 ;
  assign n9937 = n9935 | n9936 ;
  assign n10453 = n10450 & n10451 ;
  assign n10454 = n10449 | n10453 ;
  assign n10455 = n9937 | n10454 ;
  assign n10456 = n9937 & n10454 ;
  assign n32066 = ~n10456 ;
  assign n10457 = n10455 & n32066 ;
  assign n9778 = n9767 & n9776 ;
  assign n9787 = n9778 | n9786 ;
  assign n5333 = n784 & n5302 ;
  assign n5294 = x[116] & n5240 ;
  assign n6260 = x[117] & n6179 ;
  assign n9788 = n5294 | n6260 ;
  assign n9789 = x[118] & n5238 ;
  assign n9790 = n9788 | n9789 ;
  assign n9791 = n5333 | n9790 ;
  assign n32067 = ~n9791 ;
  assign n9792 = x[23] & n32067 ;
  assign n9793 = n28221 & n9791 ;
  assign n9794 = n9792 | n9793 ;
  assign n32068 = ~n9794 ;
  assign n9795 = n9787 & n32068 ;
  assign n32069 = ~n9787 ;
  assign n9797 = n32069 & n9794 ;
  assign n9798 = n9795 | n9797 ;
  assign n4479 = n452 & n4474 ;
  assign n358 = x[113] & n330 ;
  assign n428 = x[114] & n390 ;
  assign n8805 = n358 | n428 ;
  assign n8806 = x[115] & n322 ;
  assign n8807 = n8805 | n8806 ;
  assign n8808 = n4479 | n8807 ;
  assign n32070 = ~n8808 ;
  assign n8809 = x[26] & n32070 ;
  assign n8810 = n28342 & n8808 ;
  assign n8811 = n8809 | n8810 ;
  assign n9236 = n9225 & n9234 ;
  assign n9241 = n9236 | n9240 ;
  assign n9242 = n8811 | n9241 ;
  assign n9243 = n8811 & n9241 ;
  assign n32071 = ~n9243 ;
  assign n9244 = n9242 & n32071 ;
  assign n8569 = n8205 & n8567 ;
  assign n8576 = n8569 | n8575 ;
  assign n4652 = n4442 & n4632 ;
  assign n4542 = x[110] & n4514 ;
  assign n4607 = x[111] & n4572 ;
  assign n8577 = n4542 | n4607 ;
  assign n8578 = x[112] & n4504 ;
  assign n8579 = n8577 | n8578 ;
  assign n8580 = n4652 | n8579 ;
  assign n32072 = ~n8580 ;
  assign n8581 = x[29] & n32072 ;
  assign n8582 = n28483 & n8580 ;
  assign n8583 = n8581 | n8582 ;
  assign n8584 = n8576 | n8583 ;
  assign n8585 = n8576 & n8583 ;
  assign n32073 = ~n8585 ;
  assign n8586 = n8584 & n32073 ;
  assign n7562 = n7558 & n7560 ;
  assign n7573 = n7569 & n7571 ;
  assign n7574 = n7562 | n7573 ;
  assign n7005 = n6996 & n7003 ;
  assign n7006 = n6995 | n7005 ;
  assign n6614 = n6341 & n6612 ;
  assign n6625 = n6621 & n6623 ;
  assign n6626 = n6614 | n6625 ;
  assign n6085 = n6076 & n6083 ;
  assign n6086 = n6075 | n6085 ;
  assign n4876 = n4872 & n4874 ;
  assign n4887 = n4878 & n4885 ;
  assign n4888 = n4876 | n4887 ;
  assign n3337 = n3333 & n3335 ;
  assign n3348 = n3337 | n3347 ;
  assign n1724 = n1690 & n1720 ;
  assign n1583 = x[86] & n1551 ;
  assign n1661 = x[87] & n1616 ;
  assign n3255 = n1583 | n1661 ;
  assign n3256 = x[88] & n1547 ;
  assign n3257 = n3255 | n3256 ;
  assign n3258 = n1724 | n3257 ;
  assign n32074 = ~n3258 ;
  assign n3259 = x[53] & n32074 ;
  assign n3260 = n30125 & n3258 ;
  assign n3261 = n3259 | n3260 ;
  assign n1757 = n32001 & n1755 ;
  assign n1795 = n1757 | n1794 ;
  assign n922 = x[77] & n900 ;
  assign n986 = x[78] & n949 ;
  assign n1735 = n922 | n986 ;
  assign n1736 = x[79] & n881 ;
  assign n1737 = n1735 | n1736 ;
  assign n1745 = n1006 & n1741 ;
  assign n1748 = n1737 | n1745 ;
  assign n32075 = ~n1748 ;
  assign n1749 = x[62] & n32075 ;
  assign n1750 = n30886 & n1748 ;
  assign n1751 = n1749 | n1750 ;
  assign n27677 = x[75] & n27215 ;
  assign n837 = x[76] & n805 ;
  assign n1252 = n27677 | n837 ;
  assign n1254 = x[11] | n1253 ;
  assign n1255 = x[11] & n1253 ;
  assign n32076 = ~n1255 ;
  assign n1256 = n1254 & n32076 ;
  assign n32077 = ~n1252 ;
  assign n1257 = n32077 & n1256 ;
  assign n32078 = ~n1256 ;
  assign n1258 = n1252 & n32078 ;
  assign n1752 = n1257 | n1258 ;
  assign n1753 = n1751 | n1752 ;
  assign n1796 = n1751 & n1752 ;
  assign n32079 = ~n1796 ;
  assign n1797 = n1753 & n32079 ;
  assign n1798 = n1795 & n1797 ;
  assign n2064 = n1795 | n1797 ;
  assign n32080 = ~n1798 ;
  assign n2065 = n32080 & n2064 ;
  assign n1221 = n1003 & n1217 ;
  assign n1096 = x[80] & n1079 ;
  assign n1153 = x[81] & n1144 ;
  assign n2066 = n1096 | n1153 ;
  assign n2067 = x[82] & n1075 ;
  assign n2068 = n2066 | n2067 ;
  assign n2069 = n1221 | n2068 ;
  assign n32081 = ~n2069 ;
  assign n2070 = x[59] & n32081 ;
  assign n2071 = n30638 & n2069 ;
  assign n2072 = n2070 | n2071 ;
  assign n2073 = n2065 | n2072 ;
  assign n2075 = n2065 & n2072 ;
  assign n32082 = ~n2075 ;
  assign n2076 = n2073 & n32082 ;
  assign n2108 = n2097 | n2107 ;
  assign n2109 = n2076 | n2108 ;
  assign n2688 = n2076 & n2108 ;
  assign n32083 = ~n2688 ;
  assign n2689 = n2109 & n32083 ;
  assign n1462 = n1239 & n1457 ;
  assign n1377 = x[83] & n1319 ;
  assign n1413 = x[84] & n1384 ;
  assign n2690 = n1377 | n1413 ;
  assign n2691 = x[85] & n1315 ;
  assign n2692 = n2690 | n2691 ;
  assign n2693 = n1462 | n2692 ;
  assign n32084 = ~n2693 ;
  assign n2694 = x[56] & n32084 ;
  assign n2695 = n30379 & n2693 ;
  assign n2696 = n2694 | n2695 ;
  assign n2697 = n2689 | n2696 ;
  assign n2699 = n2689 & n2696 ;
  assign n32085 = ~n2699 ;
  assign n2700 = n2697 & n32085 ;
  assign n2794 = n2785 & n2792 ;
  assign n32086 = ~n2794 ;
  assign n2795 = n2784 & n32086 ;
  assign n32087 = ~n2700 ;
  assign n2796 = n32087 & n2795 ;
  assign n32088 = ~n2795 ;
  assign n3262 = n2700 & n32088 ;
  assign n3263 = n2796 | n3262 ;
  assign n32089 = ~n3261 ;
  assign n3264 = n32089 & n3263 ;
  assign n32090 = ~n3263 ;
  assign n3349 = n3261 & n32090 ;
  assign n3350 = n3264 | n3349 ;
  assign n3351 = n3348 | n3350 ;
  assign n3352 = n3348 & n3350 ;
  assign n32091 = ~n3352 ;
  assign n3669 = n3351 & n32091 ;
  assign n2051 = n2007 & n2046 ;
  assign n1909 = x[89] & n1866 ;
  assign n1969 = x[90] & n1931 ;
  assign n3670 = n1909 | n1969 ;
  assign n3671 = x[91] & n1862 ;
  assign n3672 = n3670 | n3671 ;
  assign n3673 = n2051 | n3672 ;
  assign n32092 = ~n3673 ;
  assign n3674 = x[50] & n32092 ;
  assign n3675 = n29865 & n3673 ;
  assign n3676 = n3674 | n3675 ;
  assign n3677 = n3669 | n3676 ;
  assign n3678 = n3669 & n3676 ;
  assign n32093 = ~n3678 ;
  assign n3679 = n3677 & n32093 ;
  assign n3812 = n3802 | n3811 ;
  assign n3813 = n3679 | n3812 ;
  assign n3814 = n3679 & n3812 ;
  assign n32094 = ~n3814 ;
  assign n4744 = n3813 & n32094 ;
  assign n2415 = n2321 & n2410 ;
  assign n2199 = x[92] & n2179 ;
  assign n2288 = x[93] & n2244 ;
  assign n4745 = n2199 | n2288 ;
  assign n4746 = x[94] & n2175 ;
  assign n4747 = n4745 | n4746 ;
  assign n4748 = n2415 | n4747 ;
  assign n32095 = ~n4748 ;
  assign n4749 = x[47] & n32095 ;
  assign n4750 = n29621 & n4748 ;
  assign n4751 = n4749 | n4750 ;
  assign n4752 = n4744 & n4751 ;
  assign n4889 = n4744 | n4751 ;
  assign n32096 = ~n4752 ;
  assign n5919 = n32096 & n4889 ;
  assign n32097 = ~n5919 ;
  assign n5920 = n4888 & n32097 ;
  assign n4890 = n4888 & n4889 ;
  assign n4891 = n4752 | n4890 ;
  assign n32098 = ~n4891 ;
  assign n5921 = n4889 & n32098 ;
  assign n5922 = n5920 | n5921 ;
  assign n2643 = n2438 & n2635 ;
  assign n2523 = x[95] & n2492 ;
  assign n2592 = x[96] & n2557 ;
  assign n5923 = n2523 | n2592 ;
  assign n5924 = x[97] & n2488 ;
  assign n5925 = n5923 | n5924 ;
  assign n5926 = n2643 | n5925 ;
  assign n32099 = ~n5926 ;
  assign n5927 = x[44] & n32099 ;
  assign n5928 = n29400 & n5926 ;
  assign n5929 = n5927 | n5928 ;
  assign n32100 = ~n5929 ;
  assign n5930 = n5922 & n32100 ;
  assign n32101 = ~n5922 ;
  assign n6087 = n32101 & n5929 ;
  assign n6088 = n5930 | n6087 ;
  assign n6089 = n6086 | n6088 ;
  assign n6090 = n6086 & n6088 ;
  assign n32102 = ~n6090 ;
  assign n6330 = n6089 & n32102 ;
  assign n3180 = n2466 & n3162 ;
  assign n3073 = x[98] & n3031 ;
  assign n3135 = x[99] & n3096 ;
  assign n6331 = n3073 | n3135 ;
  assign n6332 = x[100] & n3027 ;
  assign n6333 = n6331 | n6332 ;
  assign n6334 = n3180 | n6333 ;
  assign n32103 = ~n6334 ;
  assign n6335 = x[41] & n32103 ;
  assign n6336 = n29184 & n6334 ;
  assign n6337 = n6335 | n6336 ;
  assign n6338 = n6330 | n6337 ;
  assign n6339 = n6330 & n6337 ;
  assign n32104 = ~n6339 ;
  assign n6627 = n6338 & n32104 ;
  assign n32105 = ~n6626 ;
  assign n6628 = n32105 & n6627 ;
  assign n32106 = ~n6627 ;
  assign n6757 = n6626 & n32106 ;
  assign n6758 = n6628 | n6757 ;
  assign n3587 = n2626 & n3574 ;
  assign n3479 = x[101] & n3443 ;
  assign n3543 = x[102] & n3508 ;
  assign n6759 = n3479 | n3543 ;
  assign n6760 = x[103] & n3439 ;
  assign n6761 = n6759 | n6760 ;
  assign n6762 = n3587 | n6761 ;
  assign n32107 = ~n6762 ;
  assign n6763 = x[38] & n32107 ;
  assign n6764 = n28996 & n6762 ;
  assign n6765 = n6763 | n6764 ;
  assign n32108 = ~n6765 ;
  assign n6766 = n6758 & n32108 ;
  assign n32109 = ~n6758 ;
  assign n7007 = n32109 & n6765 ;
  assign n7008 = n6766 | n7007 ;
  assign n7009 = n7006 | n7008 ;
  assign n7010 = n7006 & n7008 ;
  assign n32110 = ~n7010 ;
  assign n7268 = n7009 & n32110 ;
  assign n4056 = n3223 & n4041 ;
  assign n3936 = x[104] & n3910 ;
  assign n4002 = x[105] & n3975 ;
  assign n7269 = n3936 | n4002 ;
  assign n7270 = x[106] & n3906 ;
  assign n7271 = n7269 | n7270 ;
  assign n7272 = n4056 | n7271 ;
  assign n32111 = ~n7272 ;
  assign n7273 = x[35] & n32111 ;
  assign n7274 = n28822 & n7272 ;
  assign n7275 = n7273 | n7274 ;
  assign n7276 = n7268 | n7275 ;
  assign n7575 = n7268 & n7275 ;
  assign n32112 = ~n7575 ;
  assign n7576 = n7276 & n32112 ;
  assign n32113 = ~n7574 ;
  assign n7577 = n32113 & n7576 ;
  assign n32114 = ~n7576 ;
  assign n8111 = n7574 & n32114 ;
  assign n8112 = n7577 | n8111 ;
  assign n8100 = n8096 & n8098 ;
  assign n8101 = n8095 | n8100 ;
  assign n3643 = n779 & n3639 ;
  assign n704 = x[107] & n663 ;
  assign n755 = x[108] & n720 ;
  assign n8102 = n704 | n755 ;
  assign n8103 = x[109] & n652 ;
  assign n8104 = n8102 | n8103 ;
  assign n8105 = n3643 | n8104 ;
  assign n32115 = ~n8105 ;
  assign n8106 = x[32] & n32115 ;
  assign n8107 = n28658 & n8105 ;
  assign n8108 = n8106 | n8107 ;
  assign n8109 = n8101 | n8108 ;
  assign n8110 = n8101 & n8108 ;
  assign n32116 = ~n8110 ;
  assign n8113 = n8109 & n32116 ;
  assign n8114 = n8112 & n8113 ;
  assign n8587 = n8112 | n8113 ;
  assign n8588 = n8586 & n8587 ;
  assign n32117 = ~n8114 ;
  assign n8589 = n32117 & n8588 ;
  assign n32118 = ~n8589 ;
  assign n9246 = n8586 & n32118 ;
  assign n9245 = n8587 & n32118 ;
  assign n9247 = n32117 & n9245 ;
  assign n9248 = n9246 | n9247 ;
  assign n9249 = n9244 & n9248 ;
  assign n9799 = n9244 | n9248 ;
  assign n9800 = n9798 & n9799 ;
  assign n32119 = ~n9249 ;
  assign n9801 = n32119 & n9800 ;
  assign n32120 = ~n9801 ;
  assign n10459 = n9798 & n32120 ;
  assign n10458 = n9799 & n32120 ;
  assign n10460 = n32119 & n10458 ;
  assign n10461 = n10459 | n10460 ;
  assign n10462 = n10457 & n10461 ;
  assign n11228 = n10457 | n10461 ;
  assign n11229 = n11227 & n11228 ;
  assign n32121 = ~n10462 ;
  assign n11230 = n32121 & n11229 ;
  assign n32122 = ~n11230 ;
  assign n11940 = n11227 & n32122 ;
  assign n11939 = n32121 & n11227 ;
  assign n32123 = ~n11939 ;
  assign n11941 = n11228 & n32123 ;
  assign n11942 = n32121 & n11941 ;
  assign n11943 = n11940 | n11942 ;
  assign n32124 = ~n11943 ;
  assign n11944 = n11938 & n32124 ;
  assign n32125 = ~n11938 ;
  assign n12773 = n32125 & n11943 ;
  assign n12774 = n11944 | n12773 ;
  assign n12775 = n12772 | n12774 ;
  assign n12776 = n12772 & n12774 ;
  assign n32126 = ~n12776 ;
  assign n23148 = n12775 & n32126 ;
  assign n23149 = n23147 & n23148 ;
  assign n32127 = ~n12774 ;
  assign n27753 = n12772 & n32127 ;
  assign n32128 = ~n12772 ;
  assign n27754 = n32128 & n12774 ;
  assign n27755 = n23147 | n27754 ;
  assign n27756 = n27753 | n27755 ;
  assign n32129 = ~n23149 ;
  assign n204 = n32129 & n27756 ;
  assign n23150 = n12776 | n23149 ;
  assign n11945 = n11938 & n11943 ;
  assign n11946 = n11937 | n11945 ;
  assign n8728 = n642 & n8706 ;
  assign n8675 = x[123] & n8645 ;
  assign n9858 = x[124] & n9278 ;
  assign n9924 = n8675 | n9858 ;
  assign n9925 = x[125] & n8643 ;
  assign n9926 = n9924 | n9925 ;
  assign n9927 = n8728 | n9926 ;
  assign n9928 = x[17] | n9927 ;
  assign n9929 = x[17] & n9927 ;
  assign n32130 = ~n9929 ;
  assign n9930 = n9928 & n32130 ;
  assign n10463 = n10456 | n10462 ;
  assign n32131 = ~n10463 ;
  assign n10464 = n9930 & n32131 ;
  assign n32132 = ~n9930 ;
  assign n10466 = n32132 & n10463 ;
  assign n10467 = n10464 | n10466 ;
  assign n5329 = n5047 & n5302 ;
  assign n5254 = x[117] & n5240 ;
  assign n6247 = x[118] & n6179 ;
  assign n8798 = n5254 | n6247 ;
  assign n8799 = x[119] & n5238 ;
  assign n8800 = n8798 | n8799 ;
  assign n8801 = n5329 | n8800 ;
  assign n32133 = ~n8801 ;
  assign n8802 = x[23] & n32133 ;
  assign n8803 = n28221 & n8801 ;
  assign n8804 = n8802 | n8803 ;
  assign n9250 = n9243 | n9249 ;
  assign n9251 = n8804 | n9250 ;
  assign n9252 = n8804 & n9250 ;
  assign n32134 = ~n9252 ;
  assign n9253 = n9251 & n32134 ;
  assign n4653 = n4087 & n4632 ;
  assign n4550 = x[111] & n4514 ;
  assign n4589 = x[112] & n4572 ;
  assign n7752 = n4550 | n4589 ;
  assign n7753 = x[113] & n4504 ;
  assign n7754 = n7752 | n7753 ;
  assign n7755 = n4653 | n7754 ;
  assign n7756 = x[29] | n7755 ;
  assign n7757 = x[29] & n7755 ;
  assign n32135 = ~n7757 ;
  assign n7758 = n7756 & n32135 ;
  assign n8115 = n8110 | n8114 ;
  assign n32136 = ~n8115 ;
  assign n8116 = n7758 & n32136 ;
  assign n32137 = ~n7758 ;
  assign n8118 = n32137 & n8115 ;
  assign n8119 = n8116 | n8118 ;
  assign n4063 = n3199 & n4041 ;
  assign n3951 = x[105] & n3910 ;
  assign n4035 = x[106] & n3975 ;
  assign n7017 = n3951 | n4035 ;
  assign n7018 = x[107] & n3906 ;
  assign n7019 = n7017 | n7018 ;
  assign n7020 = n4063 | n7019 ;
  assign n32138 = ~n7020 ;
  assign n7021 = x[35] & n32138 ;
  assign n7022 = n28822 & n7020 ;
  assign n7023 = n7021 | n7022 ;
  assign n6767 = n6758 & n6765 ;
  assign n7011 = n6767 | n7010 ;
  assign n3588 = n3001 & n3574 ;
  assign n3487 = x[102] & n3443 ;
  assign n3535 = x[103] & n3508 ;
  assign n6635 = n3487 | n3535 ;
  assign n6636 = x[104] & n3439 ;
  assign n6637 = n6635 | n6636 ;
  assign n6638 = n3588 | n6637 ;
  assign n6639 = x[38] | n6638 ;
  assign n6640 = x[38] & n6638 ;
  assign n32139 = ~n6640 ;
  assign n6641 = n6639 & n32139 ;
  assign n6629 = n6626 & n6627 ;
  assign n6630 = n6339 | n6629 ;
  assign n3184 = n2977 & n3162 ;
  assign n3065 = x[99] & n3031 ;
  assign n3118 = x[100] & n3096 ;
  assign n6095 = n3065 | n3118 ;
  assign n6096 = x[101] & n3027 ;
  assign n6097 = n6095 | n6096 ;
  assign n6098 = n3184 | n6097 ;
  assign n6099 = x[41] | n6098 ;
  assign n6100 = x[41] & n6098 ;
  assign n32140 = ~n6100 ;
  assign n6101 = n6099 & n32140 ;
  assign n5931 = n5922 & n5929 ;
  assign n6091 = n5931 | n6090 ;
  assign n2846 = n2635 & n2841 ;
  assign n2512 = x[96] & n2492 ;
  assign n2571 = x[97] & n2557 ;
  assign n4897 = n2512 | n2571 ;
  assign n4898 = x[98] & n2488 ;
  assign n4899 = n4897 | n4898 ;
  assign n4900 = n2846 | n4899 ;
  assign n4901 = x[44] | n4900 ;
  assign n4902 = x[44] & n4900 ;
  assign n32141 = ~n4902 ;
  assign n4903 = n4901 & n32141 ;
  assign n2329 = n2152 & n2321 ;
  assign n2201 = x[93] & n2179 ;
  assign n2278 = x[94] & n2244 ;
  assign n3820 = n2201 | n2278 ;
  assign n3821 = x[95] & n2175 ;
  assign n3822 = n3820 | n3821 ;
  assign n3823 = n2329 | n3822 ;
  assign n3824 = x[47] | n3823 ;
  assign n3825 = x[47] & n3823 ;
  assign n32142 = ~n3825 ;
  assign n3826 = n3824 & n32142 ;
  assign n3815 = n3678 | n3814 ;
  assign n867 = x[77] & n805 ;
  assign n868 = x[76] & n27215 ;
  assign n869 = n867 | n868 ;
  assign n1259 = n27892 & n1253 ;
  assign n1260 = n1258 | n1259 ;
  assign n32143 = ~n1260 ;
  assign n1261 = n869 & n32143 ;
  assign n32144 = ~n869 ;
  assign n1262 = n32144 & n1260 ;
  assign n1263 = n1261 | n1262 ;
  assign n919 = x[78] & n900 ;
  assign n959 = x[79] & n949 ;
  assign n1264 = n919 | n959 ;
  assign n1265 = x[80] & n881 ;
  assign n1266 = n1264 | n1265 ;
  assign n1274 = n1006 & n1270 ;
  assign n1275 = n1266 | n1274 ;
  assign n32145 = ~n1275 ;
  assign n1276 = x[62] & n32145 ;
  assign n1277 = n30886 & n1275 ;
  assign n1278 = n1276 | n1277 ;
  assign n32146 = ~n1278 ;
  assign n1279 = n1263 & n32146 ;
  assign n32147 = ~n1263 ;
  assign n1280 = n32147 & n1278 ;
  assign n1734 = n1279 | n1280 ;
  assign n32148 = ~n1752 ;
  assign n1754 = n1751 & n32148 ;
  assign n32149 = ~n1797 ;
  assign n1799 = n1795 & n32149 ;
  assign n1800 = n1754 | n1799 ;
  assign n32150 = ~n1800 ;
  assign n1801 = n1734 & n32150 ;
  assign n32151 = ~n1734 ;
  assign n1802 = n32151 & n1800 ;
  assign n1803 = n1801 | n1802 ;
  assign n1223 = n1057 & n1217 ;
  assign n1125 = x[81] & n1079 ;
  assign n1179 = x[82] & n1144 ;
  assign n1804 = n1125 | n1179 ;
  assign n1805 = x[83] & n1075 ;
  assign n1806 = n1804 | n1805 ;
  assign n1807 = n1223 | n1806 ;
  assign n32152 = ~n1807 ;
  assign n1808 = x[59] & n32152 ;
  assign n1809 = n30638 & n1807 ;
  assign n1810 = n1808 | n1809 ;
  assign n1811 = n1803 | n1810 ;
  assign n2062 = n1803 & n1810 ;
  assign n32153 = ~n2062 ;
  assign n2063 = n1811 & n32153 ;
  assign n32154 = ~n2065 ;
  assign n2074 = n32154 & n2072 ;
  assign n32155 = ~n2076 ;
  assign n2110 = n32155 & n2108 ;
  assign n2111 = n2074 | n2110 ;
  assign n32156 = ~n2111 ;
  assign n2112 = n2063 & n32156 ;
  assign n32157 = ~n2063 ;
  assign n2113 = n32157 & n2111 ;
  assign n2114 = n2112 | n2113 ;
  assign n1463 = n1213 & n1457 ;
  assign n1349 = x[84] & n1319 ;
  assign n1417 = x[85] & n1384 ;
  assign n2115 = n1349 | n1417 ;
  assign n2116 = x[86] & n1315 ;
  assign n2117 = n2115 | n2116 ;
  assign n2118 = n1463 | n2117 ;
  assign n32158 = ~n2118 ;
  assign n2119 = x[56] & n32158 ;
  assign n2120 = n30379 & n2118 ;
  assign n2121 = n2119 | n2120 ;
  assign n2122 = n2114 | n2121 ;
  assign n2686 = n2114 & n2121 ;
  assign n32159 = ~n2686 ;
  assign n2687 = n2122 & n32159 ;
  assign n32160 = ~n2689 ;
  assign n2698 = n32160 & n2696 ;
  assign n2797 = n2700 | n2795 ;
  assign n32161 = ~n2698 ;
  assign n2798 = n32161 & n2797 ;
  assign n2799 = n2687 & n2798 ;
  assign n2800 = n2687 | n2798 ;
  assign n32162 = ~n2799 ;
  assign n2801 = n32162 & n2800 ;
  assign n1694 = n1453 & n1690 ;
  assign n1586 = x[87] & n1551 ;
  assign n1670 = x[88] & n1616 ;
  assign n2802 = n1586 | n1670 ;
  assign n2803 = x[89] & n1547 ;
  assign n2804 = n2802 | n2803 ;
  assign n2805 = n1694 | n2804 ;
  assign n32163 = ~n2805 ;
  assign n2806 = x[53] & n32163 ;
  assign n2807 = n30125 & n2805 ;
  assign n2808 = n2806 | n2807 ;
  assign n32164 = ~n2808 ;
  assign n2809 = n2801 & n32164 ;
  assign n32165 = ~n2801 ;
  assign n3253 = n32165 & n2808 ;
  assign n3254 = n2809 | n3253 ;
  assign n3265 = n3261 & n3263 ;
  assign n3353 = n3265 | n3352 ;
  assign n3354 = n3254 | n3353 ;
  assign n3355 = n3254 & n3353 ;
  assign n32166 = ~n3355 ;
  assign n3356 = n3354 & n32166 ;
  assign n2018 = n1841 & n2007 ;
  assign n1905 = x[90] & n1866 ;
  assign n1977 = x[91] & n1931 ;
  assign n3357 = n1905 | n1977 ;
  assign n3358 = x[92] & n1862 ;
  assign n3359 = n3357 | n3358 ;
  assign n3360 = n2018 | n3359 ;
  assign n32167 = ~n3360 ;
  assign n3361 = x[50] & n32167 ;
  assign n3362 = n29865 & n3360 ;
  assign n3363 = n3361 | n3362 ;
  assign n32168 = ~n3363 ;
  assign n3364 = n3356 & n32168 ;
  assign n32169 = ~n3356 ;
  assign n3816 = n32169 & n3363 ;
  assign n3817 = n3364 | n3816 ;
  assign n32170 = ~n3815 ;
  assign n3818 = n32170 & n3817 ;
  assign n32171 = ~n3817 ;
  assign n3827 = n3815 & n32171 ;
  assign n3828 = n3818 | n3827 ;
  assign n3829 = n3826 & n3828 ;
  assign n4892 = n3818 | n3826 ;
  assign n4893 = n3827 | n4892 ;
  assign n32172 = ~n3829 ;
  assign n4894 = n32172 & n4893 ;
  assign n32173 = ~n4894 ;
  assign n4895 = n4891 & n32173 ;
  assign n4904 = n32098 & n4894 ;
  assign n4905 = n4895 | n4904 ;
  assign n4906 = n4903 & n4905 ;
  assign n6092 = n4903 | n4905 ;
  assign n32174 = ~n4906 ;
  assign n6093 = n32174 & n6092 ;
  assign n32175 = ~n6093 ;
  assign n6102 = n6091 & n32175 ;
  assign n32176 = ~n6091 ;
  assign n6103 = n32176 & n6093 ;
  assign n6104 = n6102 | n6103 ;
  assign n6105 = n6101 & n6104 ;
  assign n6631 = n6101 | n6103 ;
  assign n6632 = n6102 | n6631 ;
  assign n32177 = ~n6105 ;
  assign n6633 = n32177 & n6632 ;
  assign n32178 = ~n6633 ;
  assign n6642 = n6630 & n32178 ;
  assign n32179 = ~n6630 ;
  assign n6643 = n32179 & n6633 ;
  assign n6644 = n6642 | n6643 ;
  assign n6645 = n6641 & n6644 ;
  assign n7012 = n6641 | n6643 ;
  assign n7013 = n6642 | n7012 ;
  assign n32180 = ~n6645 ;
  assign n7014 = n32180 & n7013 ;
  assign n32181 = ~n7014 ;
  assign n7015 = n7011 & n32181 ;
  assign n32182 = ~n7011 ;
  assign n7024 = n32182 & n7014 ;
  assign n7025 = n7015 | n7024 ;
  assign n32183 = ~n7023 ;
  assign n7026 = n32183 & n7025 ;
  assign n32184 = ~n7025 ;
  assign n7591 = n7023 & n32184 ;
  assign n7592 = n7026 | n7591 ;
  assign n7578 = n7574 & n7576 ;
  assign n7579 = n7575 | n7578 ;
  assign n654 = x[110] & n652 ;
  assign n7580 = x[108] & n663 ;
  assign n7581 = x[109] & n720 ;
  assign n7582 = n7580 | n7581 ;
  assign n7583 = n654 | n7582 ;
  assign n7584 = n779 & n3615 ;
  assign n7585 = n7583 | n7584 ;
  assign n7586 = n28658 & n7585 ;
  assign n32185 = ~n7585 ;
  assign n7587 = x[32] & n32185 ;
  assign n7588 = n7586 | n7587 ;
  assign n32186 = ~n7588 ;
  assign n7589 = n7579 & n32186 ;
  assign n32187 = ~n7579 ;
  assign n7593 = n32187 & n7588 ;
  assign n7594 = n7589 | n7593 ;
  assign n7595 = n7592 | n7594 ;
  assign n7596 = n7592 & n7594 ;
  assign n32188 = ~n7596 ;
  assign n8120 = n7595 & n32188 ;
  assign n8121 = n8119 | n8120 ;
  assign n8122 = n8119 & n8120 ;
  assign n32189 = ~n8122 ;
  assign n8602 = n8121 & n32189 ;
  assign n8590 = n8585 | n8589 ;
  assign n323 = x[116] & n322 ;
  assign n8591 = x[114] & n330 ;
  assign n8592 = x[115] & n390 ;
  assign n8593 = n8591 | n8592 ;
  assign n8594 = n323 | n8593 ;
  assign n8595 = n452 & n4702 ;
  assign n8596 = n8594 | n8595 ;
  assign n8597 = n28342 & n8596 ;
  assign n32190 = ~n8596 ;
  assign n8598 = x[26] & n32190 ;
  assign n8599 = n8597 | n8598 ;
  assign n32191 = ~n8599 ;
  assign n8600 = n8590 & n32191 ;
  assign n32192 = ~n8590 ;
  assign n8603 = n32192 & n8599 ;
  assign n8604 = n8600 | n8603 ;
  assign n8605 = n8602 & n8604 ;
  assign n9254 = n8602 | n8604 ;
  assign n32193 = ~n8605 ;
  assign n9255 = n32193 & n9254 ;
  assign n32194 = ~n9255 ;
  assign n9256 = n9253 & n32194 ;
  assign n32195 = ~n9253 ;
  assign n9814 = n32195 & n9255 ;
  assign n9815 = n9256 | n9814 ;
  assign n9796 = n9787 & n9794 ;
  assign n9802 = n9796 | n9801 ;
  assign n7669 = x[122] & n7098 ;
  assign n9803 = x[120] & n7100 ;
  assign n9804 = x[121] & n7647 ;
  assign n9805 = n9803 | n9804 ;
  assign n9806 = n7669 | n9805 ;
  assign n9807 = n5022 & n7162 ;
  assign n9808 = n9806 | n9807 ;
  assign n9809 = n28114 & n9808 ;
  assign n32196 = ~n9808 ;
  assign n9810 = x[20] & n32196 ;
  assign n9811 = n9809 | n9810 ;
  assign n32197 = ~n9811 ;
  assign n9812 = n9802 & n32197 ;
  assign n32198 = ~n9802 ;
  assign n9816 = n32198 & n9811 ;
  assign n9817 = n9812 | n9816 ;
  assign n32199 = ~n9817 ;
  assign n9818 = n9815 & n32199 ;
  assign n32200 = ~n9815 ;
  assign n10468 = n32200 & n9817 ;
  assign n10469 = n9818 | n10468 ;
  assign n10470 = n10467 | n10469 ;
  assign n10471 = n10467 & n10469 ;
  assign n32201 = ~n10471 ;
  assign n11242 = n10470 & n32201 ;
  assign n11231 = n11226 | n11230 ;
  assign n10587 = n6186 & n10542 ;
  assign n11233 = x[126] & n10481 ;
  assign n11234 = x[127] & n11232 ;
  assign n11235 = n11233 | n11234 ;
  assign n11236 = n10587 | n11235 ;
  assign n32202 = ~n11236 ;
  assign n11237 = x[14] & n32202 ;
  assign n11238 = n27956 & n11236 ;
  assign n11239 = n11237 | n11238 ;
  assign n32203 = ~n11239 ;
  assign n11240 = n11231 & n32203 ;
  assign n32204 = ~n11231 ;
  assign n11243 = n32204 & n11239 ;
  assign n11244 = n11240 | n11243 ;
  assign n11245 = n11242 & n11244 ;
  assign n11947 = n11242 | n11243 ;
  assign n11948 = n11240 | n11947 ;
  assign n32205 = ~n11245 ;
  assign n11949 = n32205 & n11948 ;
  assign n32206 = ~n11949 ;
  assign n11950 = n11946 & n32206 ;
  assign n32207 = ~n11946 ;
  assign n23151 = n32207 & n11949 ;
  assign n23152 = n11950 | n23151 ;
  assign n23153 = n23150 & n23152 ;
  assign n27758 = n23150 | n23151 ;
  assign n27759 = n11950 | n27758 ;
  assign n32208 = ~n23153 ;
  assign n205 = n32208 & n27759 ;
  assign n11951 = n11946 & n11949 ;
  assign n23154 = n11951 | n23153 ;
  assign n11241 = n11231 & n11239 ;
  assign n11246 = n11241 | n11245 ;
  assign n10465 = n9930 & n10463 ;
  assign n10472 = n10465 | n10471 ;
  assign n10524 = x[127] & n10481 ;
  assign n10590 = n5360 & n10542 ;
  assign n10605 = n10524 | n10590 ;
  assign n32209 = ~n10605 ;
  assign n10606 = x[14] & n32209 ;
  assign n10607 = n27956 & n10605 ;
  assign n10608 = n10606 | n10607 ;
  assign n10609 = n10472 | n10608 ;
  assign n10610 = n10472 & n10608 ;
  assign n32210 = ~n10610 ;
  assign n10611 = n10609 & n32210 ;
  assign n7166 = n5417 & n7162 ;
  assign n7142 = x[121] & n7100 ;
  assign n7718 = x[122] & n7647 ;
  assign n8791 = n7142 | n7718 ;
  assign n8792 = x[123] & n7098 ;
  assign n8793 = n8791 | n8792 ;
  assign n8794 = n7166 | n8793 ;
  assign n8795 = x[20] | n8794 ;
  assign n8796 = x[20] & n8794 ;
  assign n32211 = ~n8796 ;
  assign n8797 = n8795 & n32211 ;
  assign n9257 = n9253 & n9255 ;
  assign n9258 = n9252 | n9257 ;
  assign n32212 = ~n9258 ;
  assign n9259 = n8797 & n32212 ;
  assign n32213 = ~n8797 ;
  assign n9261 = n32213 & n9258 ;
  assign n9262 = n9259 | n9261 ;
  assign n5346 = n4678 & n5302 ;
  assign n5271 = x[118] & n5240 ;
  assign n6251 = x[119] & n6179 ;
  assign n8192 = n5271 | n6251 ;
  assign n8193 = x[120] & n5238 ;
  assign n8194 = n8192 | n8193 ;
  assign n8195 = n5346 | n8194 ;
  assign n32214 = ~n8195 ;
  assign n8196 = x[23] & n32214 ;
  assign n8197 = n28221 & n8195 ;
  assign n8198 = n8196 | n8197 ;
  assign n8601 = n8590 & n8599 ;
  assign n8606 = n8601 | n8605 ;
  assign n8607 = n8198 | n8606 ;
  assign n8608 = n8198 & n8606 ;
  assign n32215 = ~n8608 ;
  assign n8609 = n8607 & n32215 ;
  assign n798 = n452 & n797 ;
  assign n335 = x[115] & n330 ;
  assign n426 = x[116] & n390 ;
  assign n7745 = n335 | n426 ;
  assign n7746 = x[117] & n322 ;
  assign n7747 = n7745 | n7746 ;
  assign n7748 = n798 | n7747 ;
  assign n32216 = ~n7748 ;
  assign n7749 = x[26] & n32216 ;
  assign n7750 = n28342 & n7748 ;
  assign n7751 = n7749 | n7750 ;
  assign n8117 = n7758 & n8115 ;
  assign n8123 = n8117 | n8122 ;
  assign n8124 = n7751 | n8123 ;
  assign n8125 = n7751 & n8123 ;
  assign n32217 = ~n8125 ;
  assign n8126 = n8124 & n32217 ;
  assign n7016 = n7011 & n7014 ;
  assign n7027 = n7023 & n7025 ;
  assign n7028 = n7016 | n7027 ;
  assign n653 = x[111] & n652 ;
  assign n7029 = x[109] & n663 ;
  assign n7030 = x[110] & n720 ;
  assign n7031 = n7029 | n7030 ;
  assign n7032 = n653 | n7031 ;
  assign n7033 = n779 & n4246 ;
  assign n7034 = n7032 | n7033 ;
  assign n7035 = n28658 & n7034 ;
  assign n32218 = ~n7034 ;
  assign n7036 = x[32] & n32218 ;
  assign n7037 = n7035 | n7036 ;
  assign n7038 = n7028 | n7037 ;
  assign n7039 = n7028 & n7037 ;
  assign n32219 = ~n7039 ;
  assign n7040 = n7038 & n32219 ;
  assign n4062 = n3876 & n4041 ;
  assign n3967 = x[106] & n3910 ;
  assign n3999 = x[107] & n3975 ;
  assign n6651 = n3967 | n3999 ;
  assign n6652 = x[108] & n3906 ;
  assign n6653 = n6651 | n6652 ;
  assign n6654 = n4062 | n6653 ;
  assign n32220 = ~n6654 ;
  assign n6655 = x[35] & n32220 ;
  assign n6656 = n28822 & n6654 ;
  assign n6657 = n6655 | n6656 ;
  assign n6634 = n6630 & n6633 ;
  assign n6646 = n6634 | n6645 ;
  assign n3603 = n3409 & n3574 ;
  assign n3499 = x[103] & n3443 ;
  assign n3528 = x[104] & n3508 ;
  assign n6110 = n3499 | n3528 ;
  assign n6111 = x[105] & n3439 ;
  assign n6112 = n6110 | n6111 ;
  assign n6113 = n3603 | n6112 ;
  assign n32221 = ~n6113 ;
  assign n6114 = x[38] & n32221 ;
  assign n6115 = n28996 & n6113 ;
  assign n6116 = n6114 | n6115 ;
  assign n6094 = n6091 & n6093 ;
  assign n6106 = n6094 | n6105 ;
  assign n3819 = n3815 & n3817 ;
  assign n3830 = n3819 | n3829 ;
  assign n2810 = n2801 & n2808 ;
  assign n32222 = ~n2810 ;
  assign n2811 = n2800 & n32222 ;
  assign n1696 = n1482 & n1690 ;
  assign n1610 = x[88] & n1551 ;
  assign n1644 = x[89] & n1616 ;
  assign n2129 = n1610 | n1644 ;
  assign n2130 = x[90] & n1547 ;
  assign n2131 = n2129 | n2130 ;
  assign n2132 = n1696 | n2131 ;
  assign n32223 = ~n2132 ;
  assign n2133 = x[53] & n32223 ;
  assign n2134 = n30125 & n2132 ;
  assign n2135 = n2133 | n2134 ;
  assign n32224 = ~n2114 ;
  assign n2123 = n32224 & n2121 ;
  assign n2124 = n2113 | n2123 ;
  assign n1281 = n1262 | n1280 ;
  assign n27670 = x[77] & n27215 ;
  assign n847 = x[78] & n805 ;
  assign n1018 = n27670 | n847 ;
  assign n32225 = ~n1018 ;
  assign n1019 = n869 & n32225 ;
  assign n1020 = n32144 & n1018 ;
  assign n1021 = n1019 | n1020 ;
  assign n893 = x[81] & n881 ;
  assign n1022 = x[79] & n900 ;
  assign n1023 = x[80] & n949 ;
  assign n1024 = n1022 | n1023 ;
  assign n1025 = n893 | n1024 ;
  assign n1032 = n1006 & n1029 ;
  assign n1033 = n1025 | n1032 ;
  assign n1034 = n30886 & n1033 ;
  assign n32226 = ~n1033 ;
  assign n1035 = x[62] & n32226 ;
  assign n1036 = n1034 | n1035 ;
  assign n1037 = n1021 | n1036 ;
  assign n1282 = n1021 & n1036 ;
  assign n32227 = ~n1282 ;
  assign n1283 = n1037 & n32227 ;
  assign n32228 = ~n1283 ;
  assign n1284 = n1281 & n32228 ;
  assign n32229 = ~n1281 ;
  assign n1285 = n32229 & n1283 ;
  assign n1286 = n1284 | n1285 ;
  assign n1120 = x[82] & n1079 ;
  assign n1181 = x[83] & n1144 ;
  assign n1287 = n1120 | n1181 ;
  assign n1288 = x[84] & n1075 ;
  assign n1289 = n1287 | n1288 ;
  assign n1297 = n1217 & n1293 ;
  assign n1298 = n1289 | n1297 ;
  assign n32230 = ~n1298 ;
  assign n1299 = x[59] & n32230 ;
  assign n1300 = n30638 & n1298 ;
  assign n1301 = n1299 | n1300 ;
  assign n1302 = n1286 | n1301 ;
  assign n1732 = n1286 & n1301 ;
  assign n32231 = ~n1732 ;
  assign n1733 = n1302 & n32231 ;
  assign n32232 = ~n1803 ;
  assign n1812 = n32232 & n1810 ;
  assign n1813 = n1802 | n1812 ;
  assign n32233 = ~n1813 ;
  assign n1814 = n1733 & n32233 ;
  assign n32234 = ~n1733 ;
  assign n1815 = n32234 & n1813 ;
  assign n1816 = n1814 | n1815 ;
  assign n1525 = n1457 & n1522 ;
  assign n1378 = x[85] & n1319 ;
  assign n1432 = x[86] & n1384 ;
  assign n1817 = n1378 | n1432 ;
  assign n1818 = x[87] & n1315 ;
  assign n1819 = n1817 | n1818 ;
  assign n1820 = n1525 | n1819 ;
  assign n32235 = ~n1820 ;
  assign n1821 = x[56] & n32235 ;
  assign n1822 = n30379 & n1820 ;
  assign n1823 = n1821 | n1822 ;
  assign n1824 = n1816 | n1823 ;
  assign n2125 = n1816 & n1823 ;
  assign n32236 = ~n2125 ;
  assign n2126 = n1824 & n32236 ;
  assign n2127 = n2124 | n2126 ;
  assign n2136 = n2124 & n2126 ;
  assign n32237 = ~n2136 ;
  assign n2137 = n2127 & n32237 ;
  assign n2138 = n2135 | n2137 ;
  assign n2812 = n2135 & n2137 ;
  assign n32238 = ~n2812 ;
  assign n2813 = n2138 & n32238 ;
  assign n32239 = ~n2813 ;
  assign n2814 = n2811 & n32239 ;
  assign n32240 = ~n2811 ;
  assign n2816 = n32240 & n2813 ;
  assign n2817 = n2814 | n2816 ;
  assign n2016 = n1685 & n2007 ;
  assign n1904 = x[91] & n1866 ;
  assign n1940 = x[92] & n1931 ;
  assign n2818 = n1904 | n1940 ;
  assign n2819 = x[93] & n1862 ;
  assign n2820 = n2818 | n2819 ;
  assign n2821 = n2016 | n2820 ;
  assign n32241 = ~n2821 ;
  assign n2822 = x[50] & n32241 ;
  assign n2823 = n29865 & n2821 ;
  assign n2824 = n2822 | n2823 ;
  assign n32242 = ~n2824 ;
  assign n2825 = n2817 & n32242 ;
  assign n32243 = ~n2817 ;
  assign n3251 = n32243 & n2824 ;
  assign n3252 = n2825 | n3251 ;
  assign n3365 = n3356 & n3363 ;
  assign n3366 = n3355 | n3365 ;
  assign n3367 = n3252 | n3366 ;
  assign n3368 = n3252 & n3366 ;
  assign n32244 = ~n3368 ;
  assign n3369 = n3367 & n32244 ;
  assign n2323 = n2000 & n2321 ;
  assign n2203 = x[94] & n2179 ;
  assign n2268 = x[95] & n2244 ;
  assign n3370 = n2203 | n2268 ;
  assign n3371 = x[96] & n2175 ;
  assign n3372 = n3370 | n3371 ;
  assign n3373 = n2323 | n3372 ;
  assign n32245 = ~n3373 ;
  assign n3374 = x[47] & n32245 ;
  assign n3375 = n29621 & n3373 ;
  assign n3376 = n3374 | n3375 ;
  assign n32246 = ~n3376 ;
  assign n3377 = n3369 & n32246 ;
  assign n32247 = ~n3369 ;
  assign n3831 = n32247 & n3376 ;
  assign n3832 = n3377 | n3831 ;
  assign n3833 = n3830 | n3832 ;
  assign n3834 = n3830 & n3832 ;
  assign n32248 = ~n3834 ;
  assign n3835 = n3833 & n32248 ;
  assign n2639 = n2313 & n2635 ;
  assign n2524 = x[97] & n2492 ;
  assign n2593 = x[98] & n2557 ;
  assign n3836 = n2524 | n2593 ;
  assign n3837 = x[99] & n2488 ;
  assign n3838 = n3836 | n3837 ;
  assign n3839 = n2639 | n3838 ;
  assign n32249 = ~n3839 ;
  assign n3840 = x[44] & n32249 ;
  assign n3841 = n29400 & n3839 ;
  assign n3842 = n3840 | n3841 ;
  assign n32250 = ~n3842 ;
  assign n3843 = n3835 & n32250 ;
  assign n32251 = ~n3835 ;
  assign n4742 = n32251 & n3842 ;
  assign n4743 = n3843 | n4742 ;
  assign n4896 = n4891 & n4894 ;
  assign n4907 = n4896 | n4906 ;
  assign n4908 = n4743 | n4907 ;
  assign n4909 = n4743 & n4907 ;
  assign n32252 = ~n4909 ;
  assign n4910 = n4908 & n32252 ;
  assign n3173 = n2867 & n3162 ;
  assign n3061 = x[100] & n3031 ;
  assign n3125 = x[101] & n3096 ;
  assign n4911 = n3061 | n3125 ;
  assign n4912 = x[102] & n3027 ;
  assign n4913 = n4911 | n4912 ;
  assign n4914 = n3173 | n4913 ;
  assign n32253 = ~n4914 ;
  assign n4915 = x[41] & n32253 ;
  assign n4916 = n29184 & n4914 ;
  assign n4917 = n4915 | n4916 ;
  assign n32254 = ~n4917 ;
  assign n4918 = n4910 & n32254 ;
  assign n32255 = ~n4910 ;
  assign n6107 = n32255 & n4917 ;
  assign n6108 = n4918 | n6107 ;
  assign n6109 = n6106 & n6108 ;
  assign n6117 = n6106 | n6108 ;
  assign n32256 = ~n6109 ;
  assign n6118 = n32256 & n6117 ;
  assign n32257 = ~n6116 ;
  assign n6119 = n32257 & n6118 ;
  assign n32258 = ~n6118 ;
  assign n6647 = n6116 & n32258 ;
  assign n6648 = n6119 | n6647 ;
  assign n32259 = ~n6646 ;
  assign n6649 = n32259 & n6648 ;
  assign n32260 = ~n6648 ;
  assign n6658 = n6646 & n32260 ;
  assign n6659 = n6649 | n6658 ;
  assign n32261 = ~n6657 ;
  assign n6660 = n32261 & n6659 ;
  assign n32262 = ~n6659 ;
  assign n7041 = n6657 & n32262 ;
  assign n7042 = n6660 | n7041 ;
  assign n32263 = ~n7042 ;
  assign n7043 = n7040 & n32263 ;
  assign n32264 = ~n7040 ;
  assign n7609 = n32264 & n7042 ;
  assign n7610 = n7043 | n7609 ;
  assign n7590 = n7579 & n7588 ;
  assign n7597 = n7590 | n7596 ;
  assign n4506 = x[114] & n4504 ;
  assign n7598 = x[112] & n4514 ;
  assign n7599 = x[113] & n4572 ;
  assign n7600 = n7598 | n7599 ;
  assign n7601 = n4506 | n7600 ;
  assign n7602 = n4276 & n4632 ;
  assign n7603 = n7601 | n7602 ;
  assign n7604 = n28483 & n7603 ;
  assign n32265 = ~n7603 ;
  assign n7605 = x[29] & n32265 ;
  assign n7606 = n7604 | n7605 ;
  assign n7607 = n7597 | n7606 ;
  assign n7608 = n7597 & n7606 ;
  assign n32266 = ~n7608 ;
  assign n7611 = n7607 & n32266 ;
  assign n7612 = n7610 & n7611 ;
  assign n8127 = n7610 | n7611 ;
  assign n32267 = ~n7612 ;
  assign n8128 = n32267 & n8127 ;
  assign n32268 = ~n8128 ;
  assign n8129 = n8126 & n32268 ;
  assign n32269 = ~n8126 ;
  assign n8610 = n32269 & n8128 ;
  assign n8611 = n8129 | n8610 ;
  assign n8612 = n8609 & n8611 ;
  assign n9263 = n8609 | n8611 ;
  assign n9264 = n9262 & n9263 ;
  assign n32270 = ~n8612 ;
  assign n9265 = n32270 & n9264 ;
  assign n32271 = ~n9265 ;
  assign n9835 = n9262 & n32271 ;
  assign n9834 = n9263 & n32271 ;
  assign n9836 = n32270 & n9834 ;
  assign n9837 = n9835 | n9836 ;
  assign n9813 = n9802 & n9811 ;
  assign n9819 = n9815 & n9817 ;
  assign n9820 = n9813 | n9819 ;
  assign n9821 = x[126] & n8643 ;
  assign n9824 = x[124] & n8645 ;
  assign n9825 = x[125] & n9278 ;
  assign n9826 = n9824 | n9825 ;
  assign n9827 = n9821 | n9826 ;
  assign n9828 = n5388 & n8706 ;
  assign n9829 = n9827 | n9828 ;
  assign n9830 = n28039 & n9829 ;
  assign n32272 = ~n9829 ;
  assign n9831 = x[17] & n32272 ;
  assign n9832 = n9830 | n9831 ;
  assign n32273 = ~n9832 ;
  assign n9838 = n9820 & n32273 ;
  assign n32274 = ~n9820 ;
  assign n9839 = n32274 & n9832 ;
  assign n9840 = n9838 | n9839 ;
  assign n9841 = n9837 & n9840 ;
  assign n10612 = n9837 | n9839 ;
  assign n10613 = n9838 | n10612 ;
  assign n32275 = ~n9841 ;
  assign n10614 = n32275 & n10613 ;
  assign n10615 = n10611 & n10614 ;
  assign n11247 = n10611 | n10614 ;
  assign n32276 = ~n10615 ;
  assign n11248 = n32276 & n11247 ;
  assign n32277 = ~n11246 ;
  assign n11249 = n32277 & n11248 ;
  assign n32278 = ~n11248 ;
  assign n23155 = n11246 & n32278 ;
  assign n23156 = n11249 | n23155 ;
  assign n23157 = n23154 | n23156 ;
  assign n23158 = n23154 & n23156 ;
  assign n32279 = ~n23158 ;
  assign n206 = n23157 & n32279 ;
  assign n9833 = n9820 & n9832 ;
  assign n9842 = n9833 | n9841 ;
  assign n8761 = n5629 & n8706 ;
  assign n8683 = x[125] & n8645 ;
  assign n9867 = x[126] & n9278 ;
  assign n9902 = n8683 | n9867 ;
  assign n9903 = x[127] & n8643 ;
  assign n9904 = n9902 | n9903 ;
  assign n9905 = n8761 | n9904 ;
  assign n32280 = ~n9905 ;
  assign n9906 = x[17] & n32280 ;
  assign n9907 = n28039 & n9905 ;
  assign n9908 = n9906 | n9907 ;
  assign n9909 = n9842 | n9908 ;
  assign n9910 = n9842 & n9908 ;
  assign n32281 = ~n9910 ;
  assign n9911 = n9909 & n32281 ;
  assign n7196 = n5838 & n7162 ;
  assign n7125 = x[122] & n7100 ;
  assign n7711 = x[123] & n7647 ;
  assign n8784 = n7125 | n7711 ;
  assign n8785 = x[124] & n7098 ;
  assign n8786 = n8784 | n8785 ;
  assign n8787 = n7196 | n8786 ;
  assign n32282 = ~n8787 ;
  assign n8788 = x[20] & n32282 ;
  assign n8789 = n28114 & n8787 ;
  assign n8790 = n8788 | n8789 ;
  assign n9260 = n8797 & n9258 ;
  assign n9266 = n9260 | n9265 ;
  assign n32283 = ~n9266 ;
  assign n9267 = n8790 & n32283 ;
  assign n32284 = ~n8790 ;
  assign n9268 = n32284 & n9266 ;
  assign n9269 = n9267 | n9268 ;
  assign n8613 = n8608 | n8612 ;
  assign n5314 = n4985 & n5302 ;
  assign n5263 = x[119] & n5240 ;
  assign n6250 = x[120] & n6179 ;
  assign n8614 = n5263 | n6250 ;
  assign n8615 = x[121] & n5238 ;
  assign n8616 = n8614 | n8615 ;
  assign n8617 = n5314 | n8616 ;
  assign n32285 = ~n8617 ;
  assign n8618 = x[23] & n32285 ;
  assign n8619 = n28221 & n8617 ;
  assign n8620 = n8618 | n8619 ;
  assign n32286 = ~n8620 ;
  assign n8621 = n8613 & n32286 ;
  assign n32287 = ~n8613 ;
  assign n8622 = n32287 & n8620 ;
  assign n8623 = n8621 | n8622 ;
  assign n785 = n452 & n784 ;
  assign n384 = x[116] & n330 ;
  assign n411 = x[117] & n390 ;
  assign n7738 = n384 | n411 ;
  assign n7739 = x[118] & n322 ;
  assign n7740 = n7738 | n7739 ;
  assign n7741 = n785 | n7740 ;
  assign n32288 = ~n7741 ;
  assign n7742 = x[26] & n32288 ;
  assign n7743 = n28342 & n7741 ;
  assign n7744 = n7742 | n7743 ;
  assign n8130 = n8126 & n8128 ;
  assign n8131 = n8125 | n8130 ;
  assign n8132 = n7744 | n8131 ;
  assign n8133 = n7744 & n8131 ;
  assign n32289 = ~n8133 ;
  assign n8134 = n8132 & n32289 ;
  assign n4662 = n4474 & n4632 ;
  assign n4545 = x[113] & n4514 ;
  assign n4609 = x[114] & n4572 ;
  assign n7261 = n4545 | n4609 ;
  assign n7262 = x[115] & n4504 ;
  assign n7263 = n7261 | n7262 ;
  assign n7264 = n4662 | n7263 ;
  assign n32290 = ~n7264 ;
  assign n7265 = x[29] & n32290 ;
  assign n7266 = n28483 & n7264 ;
  assign n7267 = n7265 | n7266 ;
  assign n7613 = n7608 | n7612 ;
  assign n7614 = n7267 | n7613 ;
  assign n7615 = n7267 & n7613 ;
  assign n32291 = ~n7615 ;
  assign n7616 = n7614 & n32291 ;
  assign n6120 = n6116 & n6118 ;
  assign n6121 = n6109 | n6120 ;
  assign n4919 = n4910 & n4917 ;
  assign n4920 = n4909 | n4919 ;
  assign n3844 = n3835 & n3842 ;
  assign n3845 = n3834 | n3844 ;
  assign n3378 = n3369 & n3376 ;
  assign n3379 = n3368 | n3378 ;
  assign n32292 = ~n1816 ;
  assign n1825 = n32292 & n1823 ;
  assign n1826 = n1815 | n1825 ;
  assign n27664 = x[78] & n27215 ;
  assign n848 = x[79] & n805 ;
  assign n870 = n27664 | n848 ;
  assign n871 = x[14] | n870 ;
  assign n872 = x[14] & n870 ;
  assign n32293 = ~n872 ;
  assign n873 = n871 & n32293 ;
  assign n874 = n869 & n873 ;
  assign n875 = n869 | n873 ;
  assign n32294 = ~n874 ;
  assign n876 = n32294 & n875 ;
  assign n927 = x[80] & n900 ;
  assign n972 = x[81] & n949 ;
  assign n997 = n927 | n972 ;
  assign n998 = x[82] & n881 ;
  assign n999 = n997 | n998 ;
  assign n1008 = n1003 & n1006 ;
  assign n1010 = n999 | n1008 ;
  assign n32295 = ~n1010 ;
  assign n1011 = x[62] & n32295 ;
  assign n1012 = n30886 & n1010 ;
  assign n1013 = n1011 | n1012 ;
  assign n1014 = n876 | n1013 ;
  assign n1016 = n876 & n1013 ;
  assign n32296 = ~n1016 ;
  assign n1017 = n1014 & n32296 ;
  assign n32297 = ~n1021 ;
  assign n1038 = n32297 & n1036 ;
  assign n1039 = n1020 | n1038 ;
  assign n32298 = ~n1039 ;
  assign n1040 = n1017 & n32298 ;
  assign n32299 = ~n1017 ;
  assign n1041 = n32299 & n1039 ;
  assign n1232 = n1040 | n1041 ;
  assign n1118 = x[83] & n1079 ;
  assign n1200 = x[84] & n1144 ;
  assign n1233 = n1118 | n1200 ;
  assign n1234 = x[85] & n1075 ;
  assign n1235 = n1233 | n1234 ;
  assign n1243 = n1217 & n1239 ;
  assign n1244 = n1235 | n1243 ;
  assign n32300 = ~n1244 ;
  assign n1245 = x[59] & n32300 ;
  assign n1246 = n30638 & n1244 ;
  assign n1247 = n1245 | n1246 ;
  assign n1248 = n1232 | n1247 ;
  assign n1250 = n1232 & n1247 ;
  assign n32301 = ~n1250 ;
  assign n1251 = n1248 & n32301 ;
  assign n32302 = ~n1286 ;
  assign n1303 = n32302 & n1301 ;
  assign n1304 = n1284 | n1303 ;
  assign n1305 = n1251 | n1304 ;
  assign n1712 = n1251 & n1304 ;
  assign n32303 = ~n1712 ;
  assign n1713 = n1305 & n32303 ;
  assign n1365 = x[86] & n1319 ;
  assign n1423 = x[87] & n1384 ;
  assign n1714 = n1365 | n1423 ;
  assign n1715 = x[88] & n1315 ;
  assign n1716 = n1714 | n1715 ;
  assign n1726 = n1457 & n1720 ;
  assign n1727 = n1716 | n1726 ;
  assign n32304 = ~n1727 ;
  assign n1728 = x[56] & n32304 ;
  assign n1729 = n30379 & n1727 ;
  assign n1730 = n1728 | n1729 ;
  assign n32305 = ~n1713 ;
  assign n1731 = n32305 & n1730 ;
  assign n32306 = ~n1730 ;
  assign n1827 = n1713 & n32306 ;
  assign n32307 = ~n1827 ;
  assign n1828 = n1826 & n32307 ;
  assign n32308 = ~n1731 ;
  assign n2036 = n32308 & n1828 ;
  assign n32309 = ~n2036 ;
  assign n2037 = n1826 & n32309 ;
  assign n1829 = n1731 | n1828 ;
  assign n2038 = n1827 | n1829 ;
  assign n32310 = ~n2037 ;
  assign n2039 = n32310 & n2038 ;
  assign n1593 = x[89] & n1551 ;
  assign n1638 = x[90] & n1616 ;
  assign n2040 = n1593 | n1638 ;
  assign n2041 = x[91] & n1547 ;
  assign n2042 = n2040 | n2041 ;
  assign n2053 = n1690 & n2046 ;
  assign n2054 = n2042 | n2053 ;
  assign n32311 = ~n2054 ;
  assign n2055 = x[53] & n32311 ;
  assign n2056 = n30125 & n2054 ;
  assign n2057 = n2055 | n2056 ;
  assign n2058 = n2039 | n2057 ;
  assign n2060 = n2039 & n2057 ;
  assign n32312 = ~n2060 ;
  assign n2061 = n2058 & n32312 ;
  assign n32313 = ~n2126 ;
  assign n2128 = n2124 & n32313 ;
  assign n32314 = ~n2137 ;
  assign n2139 = n2135 & n32314 ;
  assign n2140 = n2128 | n2139 ;
  assign n2141 = n2061 | n2140 ;
  assign n2673 = n2061 & n2140 ;
  assign n32315 = ~n2673 ;
  assign n2674 = n2141 & n32315 ;
  assign n2417 = n2007 & n2410 ;
  assign n1907 = x[92] & n1866 ;
  assign n1947 = x[93] & n1931 ;
  assign n2675 = n1907 | n1947 ;
  assign n2676 = x[94] & n1862 ;
  assign n2677 = n2675 | n2676 ;
  assign n2678 = n2417 | n2677 ;
  assign n32316 = ~n2678 ;
  assign n2679 = x[50] & n32316 ;
  assign n2680 = n29865 & n2678 ;
  assign n2681 = n2679 | n2680 ;
  assign n2682 = n2674 | n2681 ;
  assign n2684 = n2674 & n2681 ;
  assign n32317 = ~n2684 ;
  assign n2685 = n2682 & n32317 ;
  assign n2815 = n2811 | n2813 ;
  assign n2826 = n2817 & n2824 ;
  assign n32318 = ~n2826 ;
  assign n2827 = n2815 & n32318 ;
  assign n32319 = ~n2685 ;
  assign n2828 = n32319 & n2827 ;
  assign n32320 = ~n2827 ;
  assign n3240 = n2685 & n32320 ;
  assign n3241 = n2828 | n3240 ;
  assign n2444 = n2321 & n2438 ;
  assign n2230 = x[95] & n2179 ;
  assign n2281 = x[96] & n2244 ;
  assign n3242 = n2230 | n2281 ;
  assign n3243 = x[97] & n2175 ;
  assign n3244 = n3242 | n3243 ;
  assign n3245 = n2444 | n3244 ;
  assign n32321 = ~n3245 ;
  assign n3246 = x[47] & n32321 ;
  assign n3247 = n29621 & n3245 ;
  assign n3248 = n3246 | n3247 ;
  assign n32322 = ~n3248 ;
  assign n3249 = n3241 & n32322 ;
  assign n32323 = ~n3241 ;
  assign n3380 = n32323 & n3248 ;
  assign n3381 = n3249 | n3380 ;
  assign n3382 = n3379 | n3381 ;
  assign n3383 = n3379 & n3381 ;
  assign n32324 = ~n3383 ;
  assign n3659 = n3382 & n32324 ;
  assign n2645 = n2466 & n2635 ;
  assign n2520 = x[98] & n2492 ;
  assign n2605 = x[99] & n2557 ;
  assign n3660 = n2520 | n2605 ;
  assign n3661 = x[100] & n2488 ;
  assign n3662 = n3660 | n3661 ;
  assign n3663 = n2645 | n3662 ;
  assign n32325 = ~n3663 ;
  assign n3664 = x[44] & n32325 ;
  assign n3665 = n29400 & n3663 ;
  assign n3666 = n3664 | n3665 ;
  assign n3667 = n3659 | n3666 ;
  assign n3668 = n3659 & n3666 ;
  assign n32326 = ~n3668 ;
  assign n3846 = n3667 & n32326 ;
  assign n32327 = ~n3845 ;
  assign n3847 = n32327 & n3846 ;
  assign n32328 = ~n3846 ;
  assign n4731 = n3845 & n32328 ;
  assign n4732 = n3847 | n4731 ;
  assign n3175 = n2626 & n3162 ;
  assign n3085 = x[101] & n3031 ;
  assign n3132 = x[102] & n3096 ;
  assign n4733 = n3085 | n3132 ;
  assign n4734 = x[103] & n3027 ;
  assign n4735 = n4733 | n4734 ;
  assign n4736 = n3175 | n4735 ;
  assign n32329 = ~n4736 ;
  assign n4737 = x[41] & n32329 ;
  assign n4738 = n29184 & n4736 ;
  assign n4739 = n4737 | n4738 ;
  assign n32330 = ~n4739 ;
  assign n4740 = n4732 & n32330 ;
  assign n32331 = ~n4732 ;
  assign n4921 = n32331 & n4739 ;
  assign n4922 = n4740 | n4921 ;
  assign n4923 = n4920 | n4922 ;
  assign n4924 = n4920 & n4922 ;
  assign n32332 = ~n4924 ;
  assign n5909 = n4923 & n32332 ;
  assign n3598 = n3223 & n3574 ;
  assign n3480 = x[104] & n3443 ;
  assign n3513 = x[105] & n3508 ;
  assign n5910 = n3480 | n3513 ;
  assign n5911 = x[106] & n3439 ;
  assign n5912 = n5910 | n5911 ;
  assign n5913 = n3598 | n5912 ;
  assign n32333 = ~n5913 ;
  assign n5914 = x[38] & n32333 ;
  assign n5915 = n28996 & n5913 ;
  assign n5916 = n5914 | n5915 ;
  assign n5917 = n5909 | n5916 ;
  assign n5918 = n5909 & n5916 ;
  assign n32334 = ~n5918 ;
  assign n6122 = n5917 & n32334 ;
  assign n6123 = n6121 & n6122 ;
  assign n6317 = n6121 | n6122 ;
  assign n32335 = ~n6123 ;
  assign n6318 = n32335 & n6317 ;
  assign n4057 = n3639 & n4041 ;
  assign n3948 = x[107] & n3910 ;
  assign n4007 = x[108] & n3975 ;
  assign n6319 = n3948 | n4007 ;
  assign n6320 = x[109] & n3906 ;
  assign n6321 = n6319 | n6320 ;
  assign n6322 = n4057 | n6321 ;
  assign n32336 = ~n6322 ;
  assign n6323 = x[35] & n32336 ;
  assign n6324 = n28822 & n6322 ;
  assign n6325 = n6323 | n6324 ;
  assign n32337 = ~n6325 ;
  assign n6326 = n6318 & n32337 ;
  assign n32338 = ~n6318 ;
  assign n6328 = n32338 & n6325 ;
  assign n6329 = n6326 | n6328 ;
  assign n6650 = n6646 & n6648 ;
  assign n6661 = n6657 & n6659 ;
  assign n6662 = n6650 | n6661 ;
  assign n32339 = ~n6662 ;
  assign n6663 = n6329 & n32339 ;
  assign n32340 = ~n6329 ;
  assign n7055 = n32340 & n6662 ;
  assign n7056 = n6663 | n7055 ;
  assign n7044 = n7040 & n7042 ;
  assign n7045 = n7039 | n7044 ;
  assign n4446 = n779 & n4442 ;
  assign n698 = x[110] & n663 ;
  assign n752 = x[111] & n720 ;
  assign n7046 = n698 | n752 ;
  assign n7047 = x[112] & n652 ;
  assign n7048 = n7046 | n7047 ;
  assign n7049 = n4446 | n7048 ;
  assign n32341 = ~n7049 ;
  assign n7050 = x[32] & n32341 ;
  assign n7051 = n28658 & n7049 ;
  assign n7052 = n7050 | n7051 ;
  assign n7053 = n7045 | n7052 ;
  assign n7054 = n7045 & n7052 ;
  assign n32342 = ~n7054 ;
  assign n7057 = n7053 & n32342 ;
  assign n7058 = n7056 & n7057 ;
  assign n7617 = n7056 | n7057 ;
  assign n7618 = n7616 & n7617 ;
  assign n32343 = ~n7058 ;
  assign n7619 = n32343 & n7618 ;
  assign n32344 = ~n7619 ;
  assign n7622 = n7616 & n32344 ;
  assign n8135 = n7617 & n32344 ;
  assign n8136 = n32343 & n8135 ;
  assign n8137 = n7622 | n8136 ;
  assign n8138 = n8134 & n8137 ;
  assign n8624 = n8134 | n8137 ;
  assign n8625 = n8623 & n8624 ;
  assign n32345 = ~n8138 ;
  assign n8626 = n32345 & n8625 ;
  assign n32346 = ~n8626 ;
  assign n9270 = n8623 & n32346 ;
  assign n9271 = n8624 & n32346 ;
  assign n9272 = n32345 & n9271 ;
  assign n9273 = n9270 | n9272 ;
  assign n9275 = n9269 & n9273 ;
  assign n9274 = n9269 | n9273 ;
  assign n9913 = n9274 & n9911 ;
  assign n32347 = ~n9275 ;
  assign n9914 = n32347 & n9913 ;
  assign n32348 = ~n9914 ;
  assign n9920 = n9911 & n32348 ;
  assign n9912 = n32347 & n9911 ;
  assign n32349 = ~n9912 ;
  assign n9921 = n9274 & n32349 ;
  assign n9922 = n32347 & n9921 ;
  assign n9923 = n9920 | n9922 ;
  assign n10616 = n10610 | n10615 ;
  assign n10617 = n9923 | n10616 ;
  assign n10618 = n9923 & n10616 ;
  assign n32350 = ~n10618 ;
  assign n10619 = n10617 & n32350 ;
  assign n11250 = n11246 & n11248 ;
  assign n23159 = n11250 | n23158 ;
  assign n23160 = n10619 & n23159 ;
  assign n27762 = n10619 | n23159 ;
  assign n32351 = ~n23160 ;
  assign n207 = n32351 & n27762 ;
  assign n9276 = n8790 & n9266 ;
  assign n9277 = n9275 | n9276 ;
  assign n8749 = n6186 & n8706 ;
  assign n9279 = x[126] & n8645 ;
  assign n9280 = x[127] & n9278 ;
  assign n9281 = n9279 | n9280 ;
  assign n9282 = n8749 | n9281 ;
  assign n32352 = ~n9282 ;
  assign n9283 = x[17] & n32352 ;
  assign n9284 = n28039 & n9282 ;
  assign n9285 = n9283 | n9284 ;
  assign n32353 = ~n9285 ;
  assign n9286 = n9277 & n32353 ;
  assign n32354 = ~n9277 ;
  assign n9288 = n32354 & n9285 ;
  assign n9289 = n9286 | n9288 ;
  assign n7201 = n642 & n7162 ;
  assign n7133 = x[123] & n7100 ;
  assign n7672 = x[124] & n7647 ;
  assign n8185 = n7133 | n7672 ;
  assign n8186 = x[125] & n7098 ;
  assign n8187 = n8185 | n8186 ;
  assign n8188 = n7201 | n8187 ;
  assign n32355 = ~n8188 ;
  assign n8189 = x[20] & n32355 ;
  assign n8190 = n28114 & n8188 ;
  assign n8191 = n8189 | n8190 ;
  assign n8627 = n8613 & n8620 ;
  assign n8628 = n8626 | n8627 ;
  assign n8629 = n8191 | n8628 ;
  assign n8630 = n8191 & n8628 ;
  assign n32356 = ~n8630 ;
  assign n8631 = n8629 & n32356 ;
  assign n8139 = n8133 | n8138 ;
  assign n6220 = x[122] & n5238 ;
  assign n8140 = x[120] & n5240 ;
  assign n8141 = x[121] & n6179 ;
  assign n8142 = n8140 | n8141 ;
  assign n8143 = n6220 | n8142 ;
  assign n8144 = n5022 & n5302 ;
  assign n8145 = n8143 | n8144 ;
  assign n8146 = n28221 & n8145 ;
  assign n32357 = ~n8145 ;
  assign n8147 = x[23] & n32357 ;
  assign n8148 = n8146 | n8147 ;
  assign n8149 = n8139 | n8148 ;
  assign n8150 = n8139 & n8148 ;
  assign n32358 = ~n8150 ;
  assign n8151 = n8149 & n32358 ;
  assign n5050 = n452 & n5047 ;
  assign n372 = x[117] & n330 ;
  assign n418 = x[118] & n390 ;
  assign n7254 = n372 | n418 ;
  assign n7255 = x[119] & n322 ;
  assign n7256 = n7254 | n7255 ;
  assign n7257 = n5050 | n7256 ;
  assign n32359 = ~n7257 ;
  assign n7258 = x[26] & n32359 ;
  assign n7259 = n28342 & n7257 ;
  assign n7260 = n7258 | n7259 ;
  assign n7620 = n7615 | n7619 ;
  assign n7621 = n7260 | n7620 ;
  assign n7623 = n7260 & n7620 ;
  assign n32360 = ~n7623 ;
  assign n7624 = n7621 & n32360 ;
  assign n4706 = n4632 & n4702 ;
  assign n4532 = x[114] & n4514 ;
  assign n4606 = x[115] & n4572 ;
  assign n6750 = n4532 | n4606 ;
  assign n6751 = x[116] & n4504 ;
  assign n6752 = n6750 | n6751 ;
  assign n6753 = n4706 | n6752 ;
  assign n6754 = x[29] | n6753 ;
  assign n6755 = x[29] & n6753 ;
  assign n32361 = ~n6755 ;
  assign n6756 = n6754 & n32361 ;
  assign n7059 = n7054 | n7058 ;
  assign n32362 = ~n7059 ;
  assign n7060 = n6756 & n32362 ;
  assign n32363 = ~n6756 ;
  assign n7062 = n32363 & n7059 ;
  assign n7063 = n7060 | n7062 ;
  assign n4091 = n779 & n4087 ;
  assign n671 = x[111] & n663 ;
  assign n746 = x[112] & n720 ;
  assign n6310 = n671 | n746 ;
  assign n6311 = x[113] & n652 ;
  assign n6312 = n6310 | n6311 ;
  assign n6313 = n4091 | n6312 ;
  assign n6314 = x[32] | n6313 ;
  assign n6315 = x[32] & n6313 ;
  assign n32364 = ~n6315 ;
  assign n6316 = n6314 & n32364 ;
  assign n6327 = n6318 & n6325 ;
  assign n6664 = n6329 & n6662 ;
  assign n6665 = n6327 | n6664 ;
  assign n32365 = ~n6665 ;
  assign n6666 = n6316 & n32365 ;
  assign n32366 = ~n6316 ;
  assign n6668 = n32366 & n6665 ;
  assign n6669 = n6666 | n6668 ;
  assign n3596 = n3199 & n3574 ;
  assign n3491 = x[105] & n3443 ;
  assign n3536 = x[106] & n3508 ;
  assign n4931 = n3491 | n3536 ;
  assign n4932 = x[107] & n3439 ;
  assign n4933 = n4931 | n4932 ;
  assign n4934 = n3596 | n4933 ;
  assign n32367 = ~n4934 ;
  assign n4935 = x[38] & n32367 ;
  assign n4936 = n28996 & n4934 ;
  assign n4937 = n4935 | n4936 ;
  assign n4741 = n4732 & n4739 ;
  assign n4925 = n4741 | n4924 ;
  assign n3170 = n3001 & n3162 ;
  assign n3076 = x[102] & n3031 ;
  assign n3122 = x[103] & n3096 ;
  assign n3854 = n3076 | n3122 ;
  assign n3855 = x[104] & n3027 ;
  assign n3856 = n3854 | n3855 ;
  assign n3857 = n3170 | n3856 ;
  assign n3858 = x[41] | n3857 ;
  assign n3859 = x[41] & n3857 ;
  assign n32368 = ~n3859 ;
  assign n3860 = n3858 & n32368 ;
  assign n3848 = n3845 & n3846 ;
  assign n3849 = n3668 | n3848 ;
  assign n2982 = n2635 & n2977 ;
  assign n2538 = x[99] & n2492 ;
  assign n2560 = x[100] & n2557 ;
  assign n3388 = n2538 | n2560 ;
  assign n3389 = x[101] & n2488 ;
  assign n3390 = n3388 | n3389 ;
  assign n3391 = n2982 | n3390 ;
  assign n3392 = x[44] | n3391 ;
  assign n3393 = x[44] & n3391 ;
  assign n32369 = ~n3393 ;
  assign n3394 = n3392 & n32369 ;
  assign n3250 = n3241 & n3248 ;
  assign n3384 = n3250 | n3383 ;
  assign n1884 = x[93] & n1866 ;
  assign n1973 = x[94] & n1931 ;
  assign n2146 = n1884 | n1973 ;
  assign n2147 = x[95] & n1862 ;
  assign n2148 = n2146 | n2147 ;
  assign n2157 = n2007 & n2152 ;
  assign n2160 = n2148 | n2157 ;
  assign n2161 = x[50] | n2160 ;
  assign n2162 = x[50] & n2160 ;
  assign n32370 = ~n2162 ;
  assign n2163 = n2161 & n32370 ;
  assign n32371 = ~n876 ;
  assign n1015 = n32371 & n1013 ;
  assign n1042 = n1015 | n1041 ;
  assign n27671 = x[79] & n27215 ;
  assign n843 = x[80] & n805 ;
  assign n1043 = n27671 | n843 ;
  assign n1044 = n27956 & n870 ;
  assign n32372 = ~n873 ;
  assign n1045 = n869 & n32372 ;
  assign n1046 = n1044 | n1045 ;
  assign n1047 = n1043 | n1046 ;
  assign n1048 = n1043 & n1046 ;
  assign n32373 = ~n1048 ;
  assign n1049 = n1047 & n32373 ;
  assign n891 = x[83] & n881 ;
  assign n1050 = x[81] & n900 ;
  assign n1051 = x[82] & n949 ;
  assign n1052 = n1050 | n1051 ;
  assign n1053 = n891 | n1052 ;
  assign n1060 = n1006 & n1057 ;
  assign n1061 = n1053 | n1060 ;
  assign n1062 = n30886 & n1061 ;
  assign n32374 = ~n1061 ;
  assign n1063 = x[62] & n32374 ;
  assign n1064 = n1062 | n1063 ;
  assign n1065 = n1049 | n1064 ;
  assign n1066 = n1049 & n1064 ;
  assign n32375 = ~n1066 ;
  assign n1067 = n1065 & n32375 ;
  assign n1068 = n1042 | n1067 ;
  assign n1069 = n1042 & n1067 ;
  assign n32376 = ~n1069 ;
  assign n1070 = n1068 & n32376 ;
  assign n1132 = x[84] & n1079 ;
  assign n1188 = x[85] & n1144 ;
  assign n1207 = n1132 | n1188 ;
  assign n1208 = x[86] & n1075 ;
  assign n1209 = n1207 | n1208 ;
  assign n1222 = n1213 & n1217 ;
  assign n1225 = n1209 | n1222 ;
  assign n32377 = ~n1225 ;
  assign n1226 = x[59] & n32377 ;
  assign n1227 = n30638 & n1225 ;
  assign n1228 = n1226 | n1227 ;
  assign n1229 = n1070 | n1228 ;
  assign n1230 = n1070 & n1228 ;
  assign n32378 = ~n1230 ;
  assign n1231 = n1229 & n32378 ;
  assign n32379 = ~n1232 ;
  assign n1249 = n32379 & n1247 ;
  assign n32380 = ~n1251 ;
  assign n1306 = n32380 & n1304 ;
  assign n1307 = n1249 | n1306 ;
  assign n32381 = ~n1307 ;
  assign n1308 = n1231 & n32381 ;
  assign n32382 = ~n1231 ;
  assign n1309 = n32382 & n1307 ;
  assign n1310 = n1308 | n1309 ;
  assign n1363 = x[87] & n1319 ;
  assign n1443 = x[88] & n1384 ;
  assign n1447 = n1363 | n1443 ;
  assign n1448 = x[89] & n1315 ;
  assign n1449 = n1447 | n1448 ;
  assign n1460 = n1453 & n1457 ;
  assign n1469 = n1449 | n1460 ;
  assign n32383 = ~n1469 ;
  assign n1470 = x[56] & n32383 ;
  assign n1471 = n30379 & n1469 ;
  assign n1472 = n1470 | n1471 ;
  assign n1473 = n1310 | n1472 ;
  assign n1830 = n1310 & n1472 ;
  assign n32384 = ~n1830 ;
  assign n1831 = n1473 & n32384 ;
  assign n1832 = n1829 & n1831 ;
  assign n1833 = n1829 | n1831 ;
  assign n32385 = ~n1832 ;
  assign n1834 = n32385 & n1833 ;
  assign n1594 = x[90] & n1551 ;
  assign n1668 = x[91] & n1616 ;
  assign n1835 = n1594 | n1668 ;
  assign n1836 = x[92] & n1547 ;
  assign n1837 = n1835 | n1836 ;
  assign n1846 = n1690 & n1841 ;
  assign n1847 = n1837 | n1846 ;
  assign n32386 = ~n1847 ;
  assign n1848 = x[53] & n32386 ;
  assign n1849 = n30125 & n1847 ;
  assign n1850 = n1848 | n1849 ;
  assign n1851 = n1834 | n1850 ;
  assign n2034 = n1834 & n1850 ;
  assign n32387 = ~n2034 ;
  assign n2035 = n1851 & n32387 ;
  assign n32388 = ~n2039 ;
  assign n2059 = n32388 & n2057 ;
  assign n32389 = ~n2061 ;
  assign n2142 = n32389 & n2140 ;
  assign n2143 = n2059 | n2142 ;
  assign n2144 = n2035 | n2143 ;
  assign n2164 = n2035 & n2143 ;
  assign n32390 = ~n2164 ;
  assign n2165 = n2144 & n32390 ;
  assign n32391 = ~n2165 ;
  assign n2166 = n2163 & n32391 ;
  assign n32392 = ~n2163 ;
  assign n2671 = n32392 & n2165 ;
  assign n2672 = n2166 | n2671 ;
  assign n32393 = ~n2674 ;
  assign n2683 = n32393 & n2681 ;
  assign n2829 = n2685 | n2827 ;
  assign n32394 = ~n2683 ;
  assign n2830 = n32394 & n2829 ;
  assign n32395 = ~n2672 ;
  assign n2831 = n32395 & n2830 ;
  assign n32396 = ~n2830 ;
  assign n2833 = n2672 & n32396 ;
  assign n2834 = n2831 | n2833 ;
  assign n2204 = x[96] & n2179 ;
  assign n2286 = x[97] & n2244 ;
  assign n2835 = n2204 | n2286 ;
  assign n2836 = x[98] & n2175 ;
  assign n2837 = n2835 | n2836 ;
  assign n2847 = n2321 & n2841 ;
  assign n2851 = n2837 | n2847 ;
  assign n32397 = ~n2851 ;
  assign n2852 = x[47] & n32397 ;
  assign n2853 = n29621 & n2851 ;
  assign n2854 = n2852 | n2853 ;
  assign n32398 = ~n2854 ;
  assign n2855 = n2834 & n32398 ;
  assign n32399 = ~n2834 ;
  assign n3385 = n32399 & n2854 ;
  assign n3386 = n2855 | n3385 ;
  assign n32400 = ~n3386 ;
  assign n3395 = n3384 & n32400 ;
  assign n32401 = ~n3384 ;
  assign n3396 = n32401 & n3386 ;
  assign n3397 = n3395 | n3396 ;
  assign n3398 = n3394 & n3397 ;
  assign n3850 = n3394 | n3396 ;
  assign n3851 = n3395 | n3850 ;
  assign n32402 = ~n3398 ;
  assign n3852 = n32402 & n3851 ;
  assign n32403 = ~n3852 ;
  assign n3861 = n3849 & n32403 ;
  assign n32404 = ~n3849 ;
  assign n3862 = n32404 & n3852 ;
  assign n3863 = n3861 | n3862 ;
  assign n3864 = n3860 & n3863 ;
  assign n4926 = n3860 | n3862 ;
  assign n4927 = n3861 | n4926 ;
  assign n32405 = ~n3864 ;
  assign n4928 = n32405 & n4927 ;
  assign n32406 = ~n4928 ;
  assign n4929 = n4925 & n32406 ;
  assign n32407 = ~n4925 ;
  assign n4938 = n32407 & n4928 ;
  assign n4939 = n4929 | n4938 ;
  assign n32408 = ~n4937 ;
  assign n4940 = n32408 & n4939 ;
  assign n32409 = ~n4939 ;
  assign n5907 = n4937 & n32409 ;
  assign n5908 = n4940 | n5907 ;
  assign n6124 = n5918 | n6123 ;
  assign n32410 = ~n6124 ;
  assign n6125 = n5908 & n32410 ;
  assign n32411 = ~n5908 ;
  assign n6127 = n32411 & n6124 ;
  assign n6128 = n6125 | n6127 ;
  assign n4058 = n3615 & n4041 ;
  assign n3937 = x[108] & n3910 ;
  assign n4016 = x[109] & n3975 ;
  assign n6129 = n3937 | n4016 ;
  assign n6130 = x[110] & n3906 ;
  assign n6131 = n6129 | n6130 ;
  assign n6132 = n4058 | n6131 ;
  assign n32412 = ~n6132 ;
  assign n6133 = x[35] & n32412 ;
  assign n6134 = n28822 & n6132 ;
  assign n6135 = n6133 | n6134 ;
  assign n32413 = ~n6135 ;
  assign n6136 = n6128 & n32413 ;
  assign n32414 = ~n6128 ;
  assign n6670 = n32414 & n6135 ;
  assign n6671 = n6136 | n6670 ;
  assign n6672 = n6669 & n6671 ;
  assign n7064 = n6669 | n6671 ;
  assign n7065 = n7063 & n7064 ;
  assign n32415 = ~n6672 ;
  assign n7066 = n32415 & n7065 ;
  assign n32416 = ~n7066 ;
  assign n7626 = n7063 & n32416 ;
  assign n7625 = n7064 & n32416 ;
  assign n7627 = n32415 & n7625 ;
  assign n7628 = n7626 | n7627 ;
  assign n7629 = n7624 & n7628 ;
  assign n8152 = n7624 | n7628 ;
  assign n8153 = n8151 & n8152 ;
  assign n32417 = ~n7629 ;
  assign n8154 = n32417 & n8153 ;
  assign n32418 = ~n8154 ;
  assign n8155 = n8151 & n32418 ;
  assign n8632 = n8152 & n32418 ;
  assign n8633 = n32417 & n8632 ;
  assign n8634 = n8155 | n8633 ;
  assign n8635 = n8631 & n8634 ;
  assign n9290 = n8631 | n8634 ;
  assign n9291 = n9289 & n9290 ;
  assign n32419 = ~n8635 ;
  assign n9292 = n32419 & n9291 ;
  assign n32420 = ~n9292 ;
  assign n9298 = n9289 & n32420 ;
  assign n9297 = n9290 & n32420 ;
  assign n9299 = n32419 & n9297 ;
  assign n9300 = n9298 | n9299 ;
  assign n9915 = n9910 | n9914 ;
  assign n32421 = ~n9915 ;
  assign n9916 = n9300 & n32421 ;
  assign n32422 = ~n9300 ;
  assign n9918 = n32422 & n9915 ;
  assign n9919 = n9916 | n9918 ;
  assign n23161 = n10618 | n23160 ;
  assign n23162 = n9919 | n23161 ;
  assign n23163 = n9919 & n23161 ;
  assign n32423 = ~n23163 ;
  assign n208 = n23162 & n32423 ;
  assign n9917 = n9300 & n9915 ;
  assign n23164 = n9917 | n23163 ;
  assign n9287 = n9277 & n9285 ;
  assign n9293 = n9287 | n9292 ;
  assign n8636 = n8630 | n8635 ;
  assign n8688 = x[127] & n8645 ;
  assign n8736 = n5360 & n8706 ;
  assign n8769 = n8688 | n8736 ;
  assign n32424 = ~n8769 ;
  assign n8770 = x[17] & n32424 ;
  assign n8771 = n28039 & n8769 ;
  assign n8772 = n8770 | n8771 ;
  assign n8773 = n8636 | n8772 ;
  assign n8774 = n8636 & n8772 ;
  assign n32425 = ~n8774 ;
  assign n8775 = n8773 & n32425 ;
  assign n7188 = n5388 & n7162 ;
  assign n7121 = x[124] & n7100 ;
  assign n7698 = x[125] & n7647 ;
  assign n7731 = n7121 | n7698 ;
  assign n7732 = x[126] & n7098 ;
  assign n7733 = n7731 | n7732 ;
  assign n7734 = n7188 | n7733 ;
  assign n32426 = ~n7734 ;
  assign n7735 = x[20] & n32426 ;
  assign n7736 = n28114 & n7734 ;
  assign n7737 = n7735 | n7736 ;
  assign n8156 = n8150 | n8154 ;
  assign n8157 = n7737 | n8156 ;
  assign n8158 = n7737 & n8156 ;
  assign n32427 = ~n8158 ;
  assign n8159 = n8157 & n32427 ;
  assign n5423 = n5302 & n5417 ;
  assign n5281 = x[121] & n5240 ;
  assign n6268 = x[122] & n6179 ;
  assign n7247 = n5281 | n6268 ;
  assign n7248 = x[123] & n5238 ;
  assign n7249 = n7247 | n7248 ;
  assign n7250 = n5423 | n7249 ;
  assign n32428 = ~n7250 ;
  assign n7251 = x[23] & n32428 ;
  assign n7252 = n28221 & n7250 ;
  assign n7253 = n7251 | n7252 ;
  assign n7630 = n7623 | n7629 ;
  assign n32429 = ~n7630 ;
  assign n7631 = n7253 & n32429 ;
  assign n32430 = ~n7253 ;
  assign n7633 = n32430 & n7630 ;
  assign n7634 = n7631 | n7633 ;
  assign n4685 = n452 & n4678 ;
  assign n360 = x[118] & n330 ;
  assign n424 = x[119] & n390 ;
  assign n6743 = n360 | n424 ;
  assign n6744 = x[120] & n322 ;
  assign n6745 = n6743 | n6744 ;
  assign n6746 = n4685 | n6745 ;
  assign n32431 = ~n6746 ;
  assign n6747 = x[26] & n32431 ;
  assign n6748 = n28342 & n6746 ;
  assign n6749 = n6747 | n6748 ;
  assign n7061 = n6756 & n7059 ;
  assign n7067 = n7061 | n7066 ;
  assign n7068 = n6749 | n7067 ;
  assign n7069 = n6749 & n7067 ;
  assign n32432 = ~n7069 ;
  assign n7070 = n7068 & n32432 ;
  assign n4659 = n797 & n4632 ;
  assign n4551 = x[115] & n4514 ;
  assign n4602 = x[116] & n4572 ;
  assign n6303 = n4551 | n4602 ;
  assign n6304 = x[117] & n4504 ;
  assign n6305 = n6303 | n6304 ;
  assign n6306 = n4659 | n6305 ;
  assign n32433 = ~n6306 ;
  assign n6307 = x[29] & n32433 ;
  assign n6308 = n28483 & n6306 ;
  assign n6309 = n6307 | n6308 ;
  assign n6667 = n6316 & n6665 ;
  assign n6673 = n6667 | n6672 ;
  assign n6674 = n6309 | n6673 ;
  assign n6675 = n6309 & n6673 ;
  assign n32434 = ~n6675 ;
  assign n6676 = n6674 & n32434 ;
  assign n4278 = n779 & n4276 ;
  assign n702 = x[112] & n663 ;
  assign n745 = x[113] & n720 ;
  assign n5900 = n702 | n745 ;
  assign n5901 = x[114] & n652 ;
  assign n5902 = n5900 | n5901 ;
  assign n5903 = n4278 | n5902 ;
  assign n5904 = x[32] | n5903 ;
  assign n5905 = x[32] & n5903 ;
  assign n32435 = ~n5905 ;
  assign n5906 = n5904 & n32435 ;
  assign n6126 = n5908 & n6124 ;
  assign n6137 = n6128 & n6135 ;
  assign n6138 = n6126 | n6137 ;
  assign n32436 = ~n6138 ;
  assign n6139 = n5906 & n32436 ;
  assign n32437 = ~n5906 ;
  assign n6141 = n32437 & n6138 ;
  assign n6142 = n6139 | n6141 ;
  assign n4930 = n4925 & n4928 ;
  assign n4941 = n4937 & n4939 ;
  assign n4942 = n4930 | n4941 ;
  assign n3490 = x[106] & n3443 ;
  assign n3548 = x[107] & n3508 ;
  assign n3870 = n3490 | n3548 ;
  assign n3871 = x[108] & n3439 ;
  assign n3872 = n3870 | n3871 ;
  assign n3880 = n3574 & n3876 ;
  assign n3886 = n3872 | n3880 ;
  assign n32438 = ~n3886 ;
  assign n3887 = x[38] & n32438 ;
  assign n3888 = n28996 & n3886 ;
  assign n3889 = n3887 | n3888 ;
  assign n3853 = n3849 & n3852 ;
  assign n3865 = n3853 | n3864 ;
  assign n3053 = x[103] & n3031 ;
  assign n3110 = x[104] & n3096 ;
  assign n3403 = n3053 | n3110 ;
  assign n3404 = x[105] & n3027 ;
  assign n3405 = n3403 | n3404 ;
  assign n3410 = n3162 & n3409 ;
  assign n3420 = n3405 | n3410 ;
  assign n32439 = ~n3420 ;
  assign n3421 = x[41] & n32439 ;
  assign n3422 = n29184 & n3420 ;
  assign n3423 = n3421 | n3422 ;
  assign n3387 = n3384 & n3386 ;
  assign n3399 = n3387 | n3398 ;
  assign n32440 = ~n1310 ;
  assign n1474 = n32440 & n1472 ;
  assign n1475 = n1309 | n1474 ;
  assign n1364 = x[88] & n1319 ;
  assign n1406 = x[89] & n1384 ;
  assign n1476 = n1364 | n1406 ;
  assign n1477 = x[90] & n1315 ;
  assign n1478 = n1476 | n1477 ;
  assign n1486 = n1457 & n1482 ;
  assign n1487 = n1478 | n1486 ;
  assign n32441 = ~n1487 ;
  assign n1488 = x[56] & n32441 ;
  assign n1489 = n30379 & n1487 ;
  assign n1490 = n1488 | n1489 ;
  assign n32442 = ~n1067 ;
  assign n1491 = n1042 & n32442 ;
  assign n32443 = ~n1070 ;
  assign n1492 = n32443 & n1228 ;
  assign n1493 = n1491 | n1492 ;
  assign n1296 = n1006 & n1293 ;
  assign n912 = x[82] & n900 ;
  assign n962 = x[83] & n949 ;
  assign n1496 = n912 | n962 ;
  assign n1497 = x[84] & n881 ;
  assign n1498 = n1496 | n1497 ;
  assign n1499 = n1296 | n1498 ;
  assign n32444 = ~n1499 ;
  assign n1500 = x[62] & n32444 ;
  assign n1501 = n30886 & n1499 ;
  assign n1502 = n1500 | n1501 ;
  assign n27685 = x[80] & n27215 ;
  assign n854 = x[81] & n805 ;
  assign n1494 = n27685 | n854 ;
  assign n32445 = ~n1043 ;
  assign n1495 = n32445 & n1494 ;
  assign n32446 = ~n1494 ;
  assign n1503 = n1043 & n32446 ;
  assign n1504 = n1495 | n1503 ;
  assign n1505 = n1502 & n1504 ;
  assign n32447 = ~n1495 ;
  assign n1506 = n32447 & n1502 ;
  assign n1507 = n1503 | n1506 ;
  assign n1508 = n1495 | n1507 ;
  assign n32448 = ~n1505 ;
  assign n1509 = n32448 & n1508 ;
  assign n1510 = n32445 & n1046 ;
  assign n32449 = ~n1049 ;
  assign n1511 = n32449 & n1064 ;
  assign n1512 = n1510 | n1511 ;
  assign n1513 = n1509 | n1512 ;
  assign n1514 = n1509 & n1512 ;
  assign n32450 = ~n1514 ;
  assign n1515 = n1513 & n32450 ;
  assign n1126 = x[85] & n1079 ;
  assign n1147 = x[86] & n1144 ;
  assign n1516 = n1126 | n1147 ;
  assign n1517 = x[87] & n1075 ;
  assign n1518 = n1516 | n1517 ;
  assign n1526 = n1217 & n1522 ;
  assign n1527 = n1518 | n1526 ;
  assign n32451 = ~n1527 ;
  assign n1528 = x[59] & n32451 ;
  assign n1529 = n30638 & n1527 ;
  assign n1530 = n1528 | n1529 ;
  assign n1531 = n1515 | n1530 ;
  assign n1532 = n1515 & n1530 ;
  assign n32452 = ~n1532 ;
  assign n1533 = n1531 & n32452 ;
  assign n1534 = n1493 | n1533 ;
  assign n1535 = n1493 & n1533 ;
  assign n32453 = ~n1535 ;
  assign n1536 = n1534 & n32453 ;
  assign n1537 = n1490 | n1536 ;
  assign n1538 = n1490 & n1536 ;
  assign n32454 = ~n1538 ;
  assign n1539 = n1537 & n32454 ;
  assign n1540 = n1475 | n1539 ;
  assign n1541 = n1475 & n1539 ;
  assign n32455 = ~n1541 ;
  assign n1542 = n1540 & n32455 ;
  assign n1590 = x[91] & n1551 ;
  assign n1662 = x[92] & n1616 ;
  assign n1679 = n1590 | n1662 ;
  assign n1680 = x[93] & n1547 ;
  assign n1681 = n1679 | n1680 ;
  assign n1698 = n1685 & n1690 ;
  assign n1705 = n1681 | n1698 ;
  assign n32456 = ~n1705 ;
  assign n1706 = x[53] & n32456 ;
  assign n1707 = n30125 & n1705 ;
  assign n1708 = n1706 | n1707 ;
  assign n1709 = n1542 | n1708 ;
  assign n1710 = n1542 & n1708 ;
  assign n32457 = ~n1710 ;
  assign n1711 = n1709 & n32457 ;
  assign n32458 = ~n1834 ;
  assign n1852 = n32458 & n1850 ;
  assign n32459 = ~n1831 ;
  assign n1853 = n1829 & n32459 ;
  assign n1854 = n1852 | n1853 ;
  assign n1855 = n1711 | n1854 ;
  assign n1856 = n1711 & n1854 ;
  assign n32460 = ~n1856 ;
  assign n1857 = n1855 & n32460 ;
  assign n1897 = x[94] & n1866 ;
  assign n1971 = x[95] & n1931 ;
  assign n1994 = n1897 | n1971 ;
  assign n1995 = x[96] & n1862 ;
  assign n1996 = n1994 | n1995 ;
  assign n2020 = n2000 & n2007 ;
  assign n2027 = n1996 | n2020 ;
  assign n32461 = ~n2027 ;
  assign n2028 = x[50] & n32461 ;
  assign n2029 = n29865 & n2027 ;
  assign n2030 = n2028 | n2029 ;
  assign n2031 = n1857 | n2030 ;
  assign n2032 = n1857 & n2030 ;
  assign n32462 = ~n2032 ;
  assign n2033 = n2031 & n32462 ;
  assign n32463 = ~n2035 ;
  assign n2145 = n32463 & n2143 ;
  assign n2167 = n2145 | n2166 ;
  assign n32464 = ~n2167 ;
  assign n2168 = n2033 & n32464 ;
  assign n32465 = ~n2033 ;
  assign n2169 = n32465 & n2167 ;
  assign n2170 = n2168 | n2169 ;
  assign n2200 = x[97] & n2179 ;
  assign n2297 = x[98] & n2244 ;
  assign n2307 = n2200 | n2297 ;
  assign n2308 = x[99] & n2175 ;
  assign n2309 = n2307 | n2308 ;
  assign n2336 = n2313 & n2321 ;
  assign n2345 = n2309 | n2336 ;
  assign n32466 = ~n2345 ;
  assign n2346 = x[47] & n32466 ;
  assign n2347 = n29621 & n2345 ;
  assign n2348 = n2346 | n2347 ;
  assign n2349 = n2170 | n2348 ;
  assign n2669 = n2170 & n2348 ;
  assign n32467 = ~n2669 ;
  assign n2670 = n2349 & n32467 ;
  assign n2832 = n2672 | n2830 ;
  assign n2856 = n2834 & n2854 ;
  assign n32468 = ~n2856 ;
  assign n2857 = n2832 & n32468 ;
  assign n2858 = n2670 & n2857 ;
  assign n2859 = n2670 | n2857 ;
  assign n32469 = ~n2858 ;
  assign n2860 = n32469 & n2859 ;
  assign n2534 = x[100] & n2492 ;
  assign n2608 = x[101] & n2557 ;
  assign n2861 = n2534 | n2608 ;
  assign n2862 = x[102] & n2488 ;
  assign n2863 = n2861 | n2862 ;
  assign n2871 = n2635 & n2867 ;
  assign n2876 = n2863 | n2871 ;
  assign n32470 = ~n2876 ;
  assign n2877 = x[44] & n32470 ;
  assign n2878 = n29400 & n2876 ;
  assign n2879 = n2877 | n2878 ;
  assign n32471 = ~n2879 ;
  assign n2880 = n2860 & n32471 ;
  assign n32472 = ~n2860 ;
  assign n3400 = n32472 & n2879 ;
  assign n3401 = n2880 | n3400 ;
  assign n3402 = n3399 | n3401 ;
  assign n3424 = n3399 & n3401 ;
  assign n32473 = ~n3424 ;
  assign n3425 = n3402 & n32473 ;
  assign n32474 = ~n3423 ;
  assign n3426 = n32474 & n3425 ;
  assign n32475 = ~n3425 ;
  assign n3866 = n3423 & n32475 ;
  assign n3867 = n3426 | n3866 ;
  assign n32476 = ~n3865 ;
  assign n3868 = n32476 & n3867 ;
  assign n32477 = ~n3867 ;
  assign n3890 = n3865 & n32477 ;
  assign n3891 = n3868 | n3890 ;
  assign n32478 = ~n3889 ;
  assign n3892 = n32478 & n3891 ;
  assign n32479 = ~n3891 ;
  assign n4943 = n3889 & n32479 ;
  assign n4944 = n3892 | n4943 ;
  assign n32480 = ~n4942 ;
  assign n4945 = n32480 & n4944 ;
  assign n32481 = ~n4944 ;
  assign n4947 = n4942 & n32481 ;
  assign n4948 = n4945 | n4947 ;
  assign n4248 = n4041 & n4246 ;
  assign n3946 = x[109] & n3910 ;
  assign n4024 = x[110] & n3975 ;
  assign n4949 = n3946 | n4024 ;
  assign n4950 = x[111] & n3906 ;
  assign n4951 = n4949 | n4950 ;
  assign n4952 = n4248 | n4951 ;
  assign n32482 = ~n4952 ;
  assign n4953 = x[35] & n32482 ;
  assign n4954 = n28822 & n4952 ;
  assign n4955 = n4953 | n4954 ;
  assign n32483 = ~n4955 ;
  assign n4956 = n4948 & n32483 ;
  assign n32484 = ~n4948 ;
  assign n6143 = n32484 & n4955 ;
  assign n6144 = n4956 | n6143 ;
  assign n6145 = n6142 & n6144 ;
  assign n6677 = n6142 | n6144 ;
  assign n6678 = n6676 & n6677 ;
  assign n32485 = ~n6145 ;
  assign n6679 = n32485 & n6678 ;
  assign n32486 = ~n6679 ;
  assign n7071 = n6676 & n32486 ;
  assign n7072 = n6677 & n32486 ;
  assign n7073 = n32485 & n7072 ;
  assign n7074 = n7071 | n7073 ;
  assign n7075 = n7070 & n7074 ;
  assign n7635 = n7070 | n7074 ;
  assign n7636 = n7634 & n7635 ;
  assign n32487 = ~n7075 ;
  assign n7637 = n32487 & n7636 ;
  assign n32488 = ~n7637 ;
  assign n8160 = n7634 & n32488 ;
  assign n8161 = n7635 & n32488 ;
  assign n8162 = n32487 & n8161 ;
  assign n8163 = n8160 | n8162 ;
  assign n32489 = ~n8163 ;
  assign n8164 = n8159 & n32489 ;
  assign n32490 = ~n8159 ;
  assign n8776 = n32490 & n8163 ;
  assign n8777 = n8164 | n8776 ;
  assign n32491 = ~n8775 ;
  assign n8778 = n32491 & n8777 ;
  assign n32492 = ~n8777 ;
  assign n9294 = n8775 & n32492 ;
  assign n9295 = n8778 | n9294 ;
  assign n32493 = ~n9295 ;
  assign n23165 = n9293 & n32493 ;
  assign n32494 = ~n9293 ;
  assign n23166 = n32494 & n9295 ;
  assign n23167 = n23165 | n23166 ;
  assign n23168 = n23164 & n23167 ;
  assign n27765 = n23164 | n23166 ;
  assign n27766 = n23165 | n27765 ;
  assign n32495 = ~n23168 ;
  assign n209 = n32495 & n27766 ;
  assign n9296 = n9293 & n9295 ;
  assign n23169 = n9296 | n23168 ;
  assign n8779 = n8775 & n8777 ;
  assign n8780 = n8774 | n8779 ;
  assign n8165 = n8159 & n8163 ;
  assign n8166 = n8158 | n8165 ;
  assign n7191 = n5629 & n7162 ;
  assign n7132 = x[125] & n7100 ;
  assign n7714 = x[126] & n7647 ;
  assign n8167 = n7132 | n7714 ;
  assign n8168 = x[127] & n7098 ;
  assign n8169 = n8167 | n8168 ;
  assign n8170 = n7191 | n8169 ;
  assign n32496 = ~n8170 ;
  assign n8171 = x[20] & n32496 ;
  assign n8172 = n28114 & n8170 ;
  assign n8173 = n8171 | n8172 ;
  assign n8174 = n8166 | n8173 ;
  assign n8175 = n8166 & n8173 ;
  assign n32497 = ~n8175 ;
  assign n8176 = n8174 & n32497 ;
  assign n5843 = n5302 & n5838 ;
  assign n5265 = x[122] & n5240 ;
  assign n6271 = x[123] & n6179 ;
  assign n7240 = n5265 | n6271 ;
  assign n7241 = x[124] & n5238 ;
  assign n7242 = n7240 | n7241 ;
  assign n7243 = n5843 | n7242 ;
  assign n32498 = ~n7243 ;
  assign n7244 = x[23] & n32498 ;
  assign n7245 = n28221 & n7243 ;
  assign n7246 = n7244 | n7245 ;
  assign n7632 = n7253 & n7630 ;
  assign n7638 = n7632 | n7637 ;
  assign n7639 = n7246 | n7638 ;
  assign n7640 = n7246 & n7638 ;
  assign n32499 = ~n7640 ;
  assign n7641 = n7639 & n32499 ;
  assign n4658 = n784 & n4632 ;
  assign n4516 = x[116] & n4514 ;
  assign n4603 = x[117] & n4572 ;
  assign n6296 = n4516 | n4603 ;
  assign n6297 = x[118] & n4504 ;
  assign n6298 = n6296 | n6297 ;
  assign n6299 = n4658 | n6298 ;
  assign n32500 = ~n6299 ;
  assign n6300 = x[29] & n32500 ;
  assign n6301 = n28483 & n6299 ;
  assign n6302 = n6300 | n6301 ;
  assign n6680 = n6675 | n6679 ;
  assign n6681 = n6302 | n6680 ;
  assign n6682 = n6302 & n6680 ;
  assign n32501 = ~n6682 ;
  assign n6683 = n6681 & n32501 ;
  assign n3427 = n3423 & n3425 ;
  assign n3428 = n3424 | n3427 ;
  assign n2881 = n2860 & n2879 ;
  assign n32502 = ~n2881 ;
  assign n2882 = n2859 & n32502 ;
  assign n32503 = ~n2170 ;
  assign n2350 = n32503 & n2348 ;
  assign n2351 = n2169 | n2350 ;
  assign n32504 = ~n1509 ;
  assign n2352 = n32504 & n1512 ;
  assign n32505 = ~n1515 ;
  assign n2353 = n32505 & n1530 ;
  assign n2354 = n2352 | n2353 ;
  assign n1241 = n1006 & n1239 ;
  assign n930 = x[83] & n900 ;
  assign n982 = x[84] & n949 ;
  assign n2355 = n930 | n982 ;
  assign n2356 = x[85] & n881 ;
  assign n2357 = n2355 | n2356 ;
  assign n2358 = n1241 | n2357 ;
  assign n2359 = x[62] | n2358 ;
  assign n2360 = x[62] & n2358 ;
  assign n32506 = ~n2360 ;
  assign n2361 = n2359 & n32506 ;
  assign n27704 = x[81] & n27215 ;
  assign n830 = x[82] & n805 ;
  assign n2362 = n27704 | n830 ;
  assign n32507 = ~n2362 ;
  assign n2363 = x[17] & n32507 ;
  assign n2364 = n28039 & n2362 ;
  assign n2365 = n2363 | n2364 ;
  assign n32508 = ~n2365 ;
  assign n2366 = n1494 & n32508 ;
  assign n2367 = n32446 & n2365 ;
  assign n2368 = n2366 | n2367 ;
  assign n32509 = ~n2368 ;
  assign n2369 = n2361 & n32509 ;
  assign n32510 = ~n2361 ;
  assign n2370 = n32510 & n2368 ;
  assign n2371 = n2369 | n2370 ;
  assign n2372 = n1507 & n2371 ;
  assign n2373 = n1507 | n2371 ;
  assign n32511 = ~n2372 ;
  assign n2374 = n32511 & n2373 ;
  assign n1725 = n1217 & n1720 ;
  assign n1115 = x[86] & n1079 ;
  assign n1186 = x[87] & n1144 ;
  assign n2375 = n1115 | n1186 ;
  assign n2376 = x[88] & n1075 ;
  assign n2377 = n2375 | n2376 ;
  assign n2378 = n1725 | n2377 ;
  assign n32512 = ~n2378 ;
  assign n2379 = x[59] & n32512 ;
  assign n2380 = n30638 & n2378 ;
  assign n2381 = n2379 | n2380 ;
  assign n32513 = ~n2381 ;
  assign n2382 = n2374 & n32513 ;
  assign n32514 = ~n2374 ;
  assign n2383 = n32514 & n2381 ;
  assign n2384 = n2382 | n2383 ;
  assign n2385 = n2354 | n2384 ;
  assign n2386 = n2354 & n2384 ;
  assign n32515 = ~n2386 ;
  assign n2387 = n2385 & n32515 ;
  assign n2052 = n1457 & n2046 ;
  assign n1352 = x[89] & n1319 ;
  assign n1415 = x[90] & n1384 ;
  assign n2388 = n1352 | n1415 ;
  assign n2389 = x[91] & n1315 ;
  assign n2390 = n2388 | n2389 ;
  assign n2391 = n2052 | n2390 ;
  assign n32516 = ~n2391 ;
  assign n2392 = x[56] & n32516 ;
  assign n2393 = n30379 & n2391 ;
  assign n2394 = n2392 | n2393 ;
  assign n2395 = n2387 | n2394 ;
  assign n2396 = n2387 & n2394 ;
  assign n32517 = ~n2396 ;
  assign n2397 = n2395 & n32517 ;
  assign n32518 = ~n1533 ;
  assign n2398 = n1493 & n32518 ;
  assign n32519 = ~n1536 ;
  assign n2399 = n1490 & n32519 ;
  assign n2400 = n2398 | n2399 ;
  assign n2401 = n2397 | n2400 ;
  assign n2402 = n2397 & n2400 ;
  assign n32520 = ~n2402 ;
  assign n2403 = n2401 & n32520 ;
  assign n1588 = x[92] & n1551 ;
  assign n1648 = x[93] & n1616 ;
  assign n2404 = n1588 | n1648 ;
  assign n2405 = x[94] & n1547 ;
  assign n2406 = n2404 | n2405 ;
  assign n2413 = n1690 & n2410 ;
  assign n2419 = n2406 | n2413 ;
  assign n32521 = ~n2419 ;
  assign n2420 = x[53] & n32521 ;
  assign n2421 = n30125 & n2419 ;
  assign n2422 = n2420 | n2421 ;
  assign n2423 = n2403 | n2422 ;
  assign n2424 = n2403 & n2422 ;
  assign n32522 = ~n2424 ;
  assign n2425 = n2423 & n32522 ;
  assign n32523 = ~n1539 ;
  assign n2426 = n1475 & n32523 ;
  assign n32524 = ~n1542 ;
  assign n2427 = n32524 & n1708 ;
  assign n2428 = n2426 | n2427 ;
  assign n2429 = n2425 | n2428 ;
  assign n2430 = n2425 & n2428 ;
  assign n32525 = ~n2430 ;
  assign n2431 = n2429 & n32525 ;
  assign n1870 = x[95] & n1866 ;
  assign n1972 = x[96] & n1931 ;
  assign n2432 = n1870 | n1972 ;
  assign n2433 = x[97] & n1862 ;
  assign n2434 = n2432 | n2433 ;
  assign n2445 = n2007 & n2438 ;
  assign n2447 = n2434 | n2445 ;
  assign n32526 = ~n2447 ;
  assign n2448 = x[50] & n32526 ;
  assign n2449 = n29865 & n2447 ;
  assign n2450 = n2448 | n2449 ;
  assign n32527 = ~n1711 ;
  assign n2451 = n32527 & n1854 ;
  assign n32528 = ~n1857 ;
  assign n2452 = n32528 & n2030 ;
  assign n2453 = n2451 | n2452 ;
  assign n2454 = n2450 | n2453 ;
  assign n2455 = n2450 & n2453 ;
  assign n32529 = ~n2455 ;
  assign n2456 = n2454 & n32529 ;
  assign n32530 = ~n2431 ;
  assign n2457 = n32530 & n2456 ;
  assign n32531 = ~n2456 ;
  assign n2458 = n2431 & n32531 ;
  assign n2459 = n2457 | n2458 ;
  assign n2217 = x[98] & n2179 ;
  assign n2273 = x[99] & n2244 ;
  assign n2460 = n2217 | n2273 ;
  assign n2461 = x[100] & n2175 ;
  assign n2462 = n2460 | n2461 ;
  assign n2471 = n2321 & n2466 ;
  assign n2474 = n2462 | n2471 ;
  assign n32532 = ~n2474 ;
  assign n2475 = x[47] & n32532 ;
  assign n2476 = n29621 & n2474 ;
  assign n2477 = n2475 | n2476 ;
  assign n32533 = ~n2477 ;
  assign n2478 = n2459 & n32533 ;
  assign n32534 = ~n2459 ;
  assign n2479 = n32534 & n2477 ;
  assign n2480 = n2478 | n2479 ;
  assign n2481 = n2351 | n2480 ;
  assign n2482 = n2351 & n2480 ;
  assign n32535 = ~n2482 ;
  assign n2483 = n2481 & n32535 ;
  assign n2540 = x[101] & n2492 ;
  assign n2610 = x[102] & n2557 ;
  assign n2620 = n2540 | n2610 ;
  assign n2621 = x[103] & n2488 ;
  assign n2622 = n2620 | n2621 ;
  assign n2647 = n2626 & n2635 ;
  assign n2663 = n2622 | n2647 ;
  assign n32536 = ~n2663 ;
  assign n2664 = x[44] & n32536 ;
  assign n2665 = n29400 & n2663 ;
  assign n2666 = n2664 | n2665 ;
  assign n2667 = n2483 | n2666 ;
  assign n2883 = n2483 & n2666 ;
  assign n32537 = ~n2883 ;
  assign n2884 = n2667 & n32537 ;
  assign n2885 = n2882 & n2884 ;
  assign n2886 = n2882 | n2884 ;
  assign n32538 = ~n2885 ;
  assign n3216 = n32538 & n2886 ;
  assign n3067 = x[104] & n3031 ;
  assign n3136 = x[105] & n3096 ;
  assign n3217 = n3067 | n3136 ;
  assign n3218 = x[106] & n3027 ;
  assign n3219 = n3217 | n3218 ;
  assign n3225 = n3162 & n3223 ;
  assign n3234 = n3219 | n3225 ;
  assign n32539 = ~n3234 ;
  assign n3235 = x[41] & n32539 ;
  assign n3236 = n29184 & n3234 ;
  assign n3237 = n3235 | n3236 ;
  assign n3238 = n3216 | n3237 ;
  assign n3239 = n3216 & n3237 ;
  assign n32540 = ~n3239 ;
  assign n3429 = n3238 & n32540 ;
  assign n3430 = n3428 & n3429 ;
  assign n3631 = n3428 | n3429 ;
  assign n32541 = ~n3430 ;
  assign n3632 = n32541 & n3631 ;
  assign n3492 = x[107] & n3443 ;
  assign n3553 = x[108] & n3508 ;
  assign n3633 = n3492 | n3553 ;
  assign n3634 = x[109] & n3439 ;
  assign n3635 = n3633 | n3634 ;
  assign n3641 = n3574 & n3639 ;
  assign n3651 = n3635 | n3641 ;
  assign n32542 = ~n3651 ;
  assign n3652 = x[38] & n32542 ;
  assign n3653 = n28996 & n3651 ;
  assign n3654 = n3652 | n3653 ;
  assign n32543 = ~n3654 ;
  assign n3655 = n3632 & n32543 ;
  assign n32544 = ~n3632 ;
  assign n3657 = n32544 & n3654 ;
  assign n3658 = n3655 | n3657 ;
  assign n3869 = n3865 & n3867 ;
  assign n3893 = n3889 & n3891 ;
  assign n3894 = n3869 | n3893 ;
  assign n32545 = ~n3894 ;
  assign n3895 = n3658 & n32545 ;
  assign n32546 = ~n3658 ;
  assign n4718 = n32546 & n3894 ;
  assign n4719 = n3895 | n4718 ;
  assign n4445 = n4041 & n4442 ;
  assign n3941 = x[110] & n3910 ;
  assign n3993 = x[111] & n3975 ;
  assign n4720 = n3941 | n3993 ;
  assign n4721 = x[112] & n3906 ;
  assign n4722 = n4720 | n4721 ;
  assign n4723 = n4445 | n4722 ;
  assign n32547 = ~n4723 ;
  assign n4724 = x[35] & n32547 ;
  assign n4725 = n28822 & n4723 ;
  assign n4726 = n4724 | n4725 ;
  assign n32548 = ~n4726 ;
  assign n4727 = n4719 & n32548 ;
  assign n32549 = ~n4719 ;
  assign n4729 = n32549 & n4726 ;
  assign n4730 = n4727 | n4729 ;
  assign n4946 = n4942 & n4944 ;
  assign n4957 = n4948 & n4955 ;
  assign n4958 = n4946 | n4957 ;
  assign n32550 = ~n4958 ;
  assign n4959 = n4730 & n32550 ;
  assign n32551 = ~n4730 ;
  assign n6149 = n32551 & n4958 ;
  assign n6150 = n4959 | n6149 ;
  assign n4480 = n779 & n4474 ;
  assign n700 = x[113] & n663 ;
  assign n741 = x[114] & n720 ;
  assign n5893 = n700 | n741 ;
  assign n5894 = x[115] & n652 ;
  assign n5895 = n5893 | n5894 ;
  assign n5896 = n4480 | n5895 ;
  assign n32552 = ~n5896 ;
  assign n5897 = x[32] & n32552 ;
  assign n5898 = n28658 & n5896 ;
  assign n5899 = n5897 | n5898 ;
  assign n6140 = n5906 & n6138 ;
  assign n6146 = n6140 | n6145 ;
  assign n6147 = n5899 | n6146 ;
  assign n6148 = n5899 & n6146 ;
  assign n32553 = ~n6148 ;
  assign n6151 = n6147 & n32553 ;
  assign n6152 = n6150 & n6151 ;
  assign n6684 = n6150 | n6151 ;
  assign n32554 = ~n6152 ;
  assign n6685 = n32554 & n6684 ;
  assign n32555 = ~n6685 ;
  assign n6686 = n6683 & n32555 ;
  assign n32556 = ~n6683 ;
  assign n7079 = n32556 & n6685 ;
  assign n7080 = n6686 | n7079 ;
  assign n4991 = n452 & n4985 ;
  assign n362 = x[119] & n330 ;
  assign n420 = x[120] & n390 ;
  assign n6736 = n362 | n420 ;
  assign n6737 = x[121] & n322 ;
  assign n6738 = n6736 | n6737 ;
  assign n6739 = n4991 | n6738 ;
  assign n32557 = ~n6739 ;
  assign n6740 = x[26] & n32557 ;
  assign n6741 = n28342 & n6739 ;
  assign n6742 = n6740 | n6741 ;
  assign n7076 = n7069 | n7075 ;
  assign n7077 = n6742 | n7076 ;
  assign n7078 = n6742 & n7076 ;
  assign n32558 = ~n7078 ;
  assign n7081 = n7077 & n32558 ;
  assign n7082 = n7080 & n7081 ;
  assign n7642 = n7080 | n7081 ;
  assign n32559 = ~n7082 ;
  assign n7643 = n32559 & n7642 ;
  assign n32560 = ~n7643 ;
  assign n7644 = n7641 & n32560 ;
  assign n32561 = ~n7641 ;
  assign n8177 = n32561 & n7643 ;
  assign n8178 = n7644 | n8177 ;
  assign n32562 = ~n8178 ;
  assign n8180 = n8176 & n32562 ;
  assign n32563 = ~n8176 ;
  assign n8781 = n32563 & n8178 ;
  assign n8782 = n8180 | n8781 ;
  assign n32564 = ~n8782 ;
  assign n23170 = n8780 & n32564 ;
  assign n32565 = ~n8780 ;
  assign n23171 = n32565 & n8782 ;
  assign n23172 = n23170 | n23171 ;
  assign n23173 = n23169 & n23172 ;
  assign n27768 = n23169 | n23171 ;
  assign n27769 = n23170 | n27768 ;
  assign n32566 = ~n23173 ;
  assign n210 = n32566 & n27769 ;
  assign n8783 = n8780 & n8782 ;
  assign n23174 = n8783 | n23173 ;
  assign n8179 = n8176 & n8178 ;
  assign n8181 = n8175 | n8179 ;
  assign n5339 = n642 & n5302 ;
  assign n5297 = x[123] & n5240 ;
  assign n6262 = x[124] & n6179 ;
  assign n6729 = n5297 | n6262 ;
  assign n6730 = x[125] & n5238 ;
  assign n6731 = n6729 | n6730 ;
  assign n6732 = n5339 | n6731 ;
  assign n32567 = ~n6732 ;
  assign n6733 = x[23] & n32567 ;
  assign n6734 = n28221 & n6732 ;
  assign n6735 = n6733 | n6734 ;
  assign n7083 = n7078 | n7082 ;
  assign n7084 = n6735 | n7083 ;
  assign n7085 = n6735 & n7083 ;
  assign n32568 = ~n7085 ;
  assign n7086 = n7084 & n32568 ;
  assign n5030 = n452 & n5022 ;
  assign n369 = x[120] & n330 ;
  assign n412 = x[121] & n390 ;
  assign n6289 = n369 | n412 ;
  assign n6290 = x[122] & n322 ;
  assign n6291 = n6289 | n6290 ;
  assign n6292 = n5030 | n6291 ;
  assign n32569 = ~n6292 ;
  assign n6293 = x[26] & n32569 ;
  assign n6294 = n28342 & n6292 ;
  assign n6295 = n6293 | n6294 ;
  assign n6687 = n6683 & n6685 ;
  assign n6688 = n6682 | n6687 ;
  assign n6689 = n6295 | n6688 ;
  assign n6690 = n6295 & n6688 ;
  assign n32570 = ~n6690 ;
  assign n6691 = n6689 & n32570 ;
  assign n5049 = n4632 & n5047 ;
  assign n4528 = x[117] & n4514 ;
  assign n4592 = x[118] & n4572 ;
  assign n5886 = n4528 | n4592 ;
  assign n5887 = x[119] & n4504 ;
  assign n5888 = n5886 | n5887 ;
  assign n5889 = n5049 | n5888 ;
  assign n5890 = x[29] | n5889 ;
  assign n5891 = x[29] & n5889 ;
  assign n32571 = ~n5891 ;
  assign n5892 = n5890 & n32571 ;
  assign n6153 = n6148 | n6152 ;
  assign n32572 = ~n6153 ;
  assign n6154 = n5892 & n32572 ;
  assign n32573 = ~n5892 ;
  assign n6156 = n32573 & n6153 ;
  assign n6157 = n6154 | n6156 ;
  assign n694 = x[114] & n663 ;
  assign n740 = x[115] & n720 ;
  assign n4696 = n694 | n740 ;
  assign n4697 = x[116] & n652 ;
  assign n4698 = n4696 | n4697 ;
  assign n4711 = n779 & n4702 ;
  assign n4714 = n4698 | n4711 ;
  assign n4715 = x[32] | n4714 ;
  assign n4716 = x[32] & n4714 ;
  assign n32574 = ~n4716 ;
  assign n4717 = n4715 & n32574 ;
  assign n4728 = n4719 & n4726 ;
  assign n4960 = n4730 & n4958 ;
  assign n4961 = n4728 | n4960 ;
  assign n32575 = ~n4961 ;
  assign n4962 = n4717 & n32575 ;
  assign n32576 = ~n4717 ;
  assign n4964 = n32576 & n4961 ;
  assign n4965 = n4962 | n4964 ;
  assign n32577 = ~n2483 ;
  assign n2668 = n32577 & n2666 ;
  assign n32578 = ~n2668 ;
  assign n2887 = n32578 & n2886 ;
  assign n2546 = x[102] & n2492 ;
  assign n2597 = x[103] & n2557 ;
  assign n2995 = n2546 | n2597 ;
  assign n2996 = x[104] & n2488 ;
  assign n2997 = n2995 | n2996 ;
  assign n3006 = n2635 & n3001 ;
  assign n3011 = n2997 | n3006 ;
  assign n3012 = x[44] | n3011 ;
  assign n3013 = x[44] & n3011 ;
  assign n32579 = ~n3013 ;
  assign n3014 = n3012 & n32579 ;
  assign n32580 = ~n2480 ;
  assign n2888 = n2351 & n32580 ;
  assign n2889 = n2479 | n2888 ;
  assign n32581 = ~n2384 ;
  assign n2890 = n2354 & n32581 ;
  assign n2891 = n2383 | n2890 ;
  assign n27720 = x[82] & n27215 ;
  assign n844 = x[83] & n805 ;
  assign n2892 = n27720 | n844 ;
  assign n2893 = n2364 | n2366 ;
  assign n32582 = ~n2893 ;
  assign n2894 = n2892 & n32582 ;
  assign n32583 = ~n2892 ;
  assign n2895 = n32583 & n2893 ;
  assign n2896 = n2894 | n2895 ;
  assign n1215 = n1006 & n1213 ;
  assign n935 = x[84] & n900 ;
  assign n979 = x[85] & n949 ;
  assign n2897 = n935 | n979 ;
  assign n2898 = x[86] & n881 ;
  assign n2899 = n2897 | n2898 ;
  assign n2900 = n1215 | n2899 ;
  assign n32584 = ~n2900 ;
  assign n2901 = x[62] & n32584 ;
  assign n2902 = n30886 & n2900 ;
  assign n2903 = n2901 | n2902 ;
  assign n2904 = n2896 | n2903 ;
  assign n2905 = n2896 & n2903 ;
  assign n32585 = ~n2905 ;
  assign n2906 = n2904 & n32585 ;
  assign n32586 = ~n2371 ;
  assign n2907 = n1507 & n32586 ;
  assign n2908 = n2369 | n2907 ;
  assign n2909 = n2906 | n2908 ;
  assign n2910 = n2906 & n2908 ;
  assign n32587 = ~n2910 ;
  assign n2911 = n2909 & n32587 ;
  assign n1455 = n1217 & n1453 ;
  assign n1081 = x[87] & n1079 ;
  assign n1173 = x[88] & n1144 ;
  assign n2912 = n1081 | n1173 ;
  assign n2913 = x[89] & n1075 ;
  assign n2914 = n2912 | n2913 ;
  assign n2915 = n1455 | n2914 ;
  assign n32588 = ~n2915 ;
  assign n2916 = x[59] & n32588 ;
  assign n2917 = n30638 & n2915 ;
  assign n2918 = n2916 | n2917 ;
  assign n2919 = n2911 | n2918 ;
  assign n2920 = n2911 & n2918 ;
  assign n32589 = ~n2920 ;
  assign n2921 = n2919 & n32589 ;
  assign n2922 = n2891 & n2921 ;
  assign n2923 = n2891 | n2921 ;
  assign n32590 = ~n2922 ;
  assign n2924 = n32590 & n2923 ;
  assign n1843 = n1457 & n1841 ;
  assign n1360 = x[90] & n1319 ;
  assign n1425 = x[91] & n1384 ;
  assign n2925 = n1360 | n1425 ;
  assign n2926 = x[92] & n1315 ;
  assign n2927 = n2925 | n2926 ;
  assign n2928 = n1843 | n2927 ;
  assign n32591 = ~n2928 ;
  assign n2929 = x[56] & n32591 ;
  assign n2930 = n30379 & n2928 ;
  assign n2931 = n2929 | n2930 ;
  assign n2932 = n2924 | n2931 ;
  assign n2933 = n2924 & n2931 ;
  assign n32592 = ~n2933 ;
  assign n2934 = n2932 & n32592 ;
  assign n32593 = ~n2387 ;
  assign n2935 = n32593 & n2394 ;
  assign n32594 = ~n2397 ;
  assign n2936 = n32594 & n2400 ;
  assign n2937 = n2935 | n2936 ;
  assign n2938 = n2934 | n2937 ;
  assign n2939 = n2934 & n2937 ;
  assign n32595 = ~n2939 ;
  assign n2940 = n2938 & n32595 ;
  assign n2156 = n1690 & n2152 ;
  assign n1585 = x[93] & n1551 ;
  assign n1665 = x[94] & n1616 ;
  assign n2941 = n1585 | n1665 ;
  assign n2942 = x[95] & n1547 ;
  assign n2943 = n2941 | n2942 ;
  assign n2944 = n2156 | n2943 ;
  assign n32596 = ~n2944 ;
  assign n2945 = x[53] & n32596 ;
  assign n2946 = n30125 & n2944 ;
  assign n2947 = n2945 | n2946 ;
  assign n2948 = n2940 | n2947 ;
  assign n2949 = n2940 & n2947 ;
  assign n32597 = ~n2949 ;
  assign n2950 = n2948 & n32597 ;
  assign n32598 = ~n2403 ;
  assign n2951 = n32598 & n2422 ;
  assign n32599 = ~n2425 ;
  assign n2952 = n32599 & n2428 ;
  assign n2953 = n2951 | n2952 ;
  assign n32600 = ~n2953 ;
  assign n2954 = n2950 & n32600 ;
  assign n32601 = ~n2950 ;
  assign n2955 = n32601 & n2953 ;
  assign n2956 = n2954 | n2955 ;
  assign n2845 = n2007 & n2841 ;
  assign n1872 = x[96] & n1866 ;
  assign n1956 = x[97] & n1931 ;
  assign n2957 = n1872 | n1956 ;
  assign n2958 = x[98] & n1862 ;
  assign n2959 = n2957 | n2958 ;
  assign n2960 = n2845 | n2959 ;
  assign n32602 = ~n2960 ;
  assign n2961 = x[50] & n32602 ;
  assign n2962 = n29865 & n2960 ;
  assign n2963 = n2961 | n2962 ;
  assign n2964 = n2956 | n2963 ;
  assign n2965 = n2956 & n2963 ;
  assign n32603 = ~n2965 ;
  assign n2966 = n2964 & n32603 ;
  assign n2967 = n2455 | n2457 ;
  assign n32604 = ~n2967 ;
  assign n2968 = n2966 & n32604 ;
  assign n32605 = ~n2966 ;
  assign n2969 = n32605 & n2967 ;
  assign n2970 = n2968 | n2969 ;
  assign n2206 = x[99] & n2179 ;
  assign n2279 = x[100] & n2244 ;
  assign n2971 = n2206 | n2279 ;
  assign n2972 = x[101] & n2175 ;
  assign n2973 = n2971 | n2972 ;
  assign n2980 = n2321 & n2977 ;
  assign n2986 = n2973 | n2980 ;
  assign n32606 = ~n2986 ;
  assign n2987 = x[47] & n32606 ;
  assign n2988 = n29621 & n2986 ;
  assign n2989 = n2987 | n2988 ;
  assign n2990 = n2970 | n2989 ;
  assign n2991 = n2970 & n2989 ;
  assign n32607 = ~n2991 ;
  assign n2992 = n2990 & n32607 ;
  assign n2993 = n2889 | n2992 ;
  assign n2994 = n2889 & n2992 ;
  assign n32608 = ~n2994 ;
  assign n3015 = n2993 & n32608 ;
  assign n32609 = ~n3015 ;
  assign n3016 = n3014 & n32609 ;
  assign n32610 = ~n3014 ;
  assign n3017 = n2993 & n32610 ;
  assign n3018 = n32608 & n3017 ;
  assign n3019 = n3016 | n3018 ;
  assign n32611 = ~n2887 ;
  assign n3020 = n32611 & n3019 ;
  assign n32612 = ~n3019 ;
  assign n3021 = n2887 & n32612 ;
  assign n3022 = n3020 | n3021 ;
  assign n3079 = x[105] & n3031 ;
  assign n3138 = x[106] & n3096 ;
  assign n3159 = n3079 | n3138 ;
  assign n3160 = x[107] & n3027 ;
  assign n3161 = n3159 | n3160 ;
  assign n3203 = n3162 & n3199 ;
  assign n3209 = n3161 | n3203 ;
  assign n32613 = ~n3209 ;
  assign n3210 = x[41] & n32613 ;
  assign n3211 = n29184 & n3209 ;
  assign n3212 = n3210 | n3211 ;
  assign n32614 = ~n3212 ;
  assign n3213 = n3022 & n32614 ;
  assign n32615 = ~n3022 ;
  assign n3214 = n32615 & n3212 ;
  assign n3215 = n3213 | n3214 ;
  assign n3431 = n3239 | n3430 ;
  assign n32616 = ~n3431 ;
  assign n3432 = n3215 & n32616 ;
  assign n32617 = ~n3215 ;
  assign n3433 = n32617 & n3431 ;
  assign n3434 = n3432 | n3433 ;
  assign n3494 = x[108] & n3443 ;
  assign n3537 = x[109] & n3508 ;
  assign n3571 = n3494 | n3537 ;
  assign n3572 = x[110] & n3439 ;
  assign n3573 = n3571 | n3572 ;
  assign n3617 = n3574 & n3615 ;
  assign n3624 = n3573 | n3617 ;
  assign n32618 = ~n3624 ;
  assign n3625 = x[38] & n32618 ;
  assign n3626 = n28996 & n3624 ;
  assign n3627 = n3625 | n3626 ;
  assign n32619 = ~n3627 ;
  assign n3628 = n3434 & n32619 ;
  assign n32620 = ~n3434 ;
  assign n3629 = n32620 & n3627 ;
  assign n3630 = n3628 | n3629 ;
  assign n3656 = n3632 & n3654 ;
  assign n3896 = n3658 & n3894 ;
  assign n3897 = n3656 | n3896 ;
  assign n32621 = ~n3897 ;
  assign n3898 = n3630 & n32621 ;
  assign n32622 = ~n3630 ;
  assign n3900 = n32622 & n3897 ;
  assign n3901 = n3898 | n3900 ;
  assign n3924 = x[111] & n3910 ;
  assign n4020 = x[112] & n3975 ;
  assign n4038 = n3924 | n4020 ;
  assign n4039 = x[113] & n3906 ;
  assign n4040 = n4038 | n4039 ;
  assign n4089 = n4041 & n4087 ;
  assign n4100 = n4040 | n4089 ;
  assign n32623 = ~n4100 ;
  assign n4101 = x[35] & n32623 ;
  assign n4102 = n28822 & n4100 ;
  assign n4103 = n4101 | n4102 ;
  assign n32624 = ~n4103 ;
  assign n4104 = n3901 & n32624 ;
  assign n32625 = ~n3901 ;
  assign n4966 = n32625 & n4103 ;
  assign n4967 = n4104 | n4966 ;
  assign n4968 = n4965 & n4967 ;
  assign n6158 = n4965 | n4967 ;
  assign n6159 = n6157 & n6158 ;
  assign n32626 = ~n4968 ;
  assign n6160 = n32626 & n6159 ;
  assign n32627 = ~n6160 ;
  assign n6692 = n6157 & n32627 ;
  assign n6693 = n6158 & n32627 ;
  assign n6694 = n32626 & n6693 ;
  assign n6695 = n6692 | n6694 ;
  assign n6696 = n6691 & n6695 ;
  assign n7087 = n6691 | n6695 ;
  assign n7088 = n7086 & n7087 ;
  assign n32628 = ~n6696 ;
  assign n7089 = n32628 & n7088 ;
  assign n32629 = ~n7089 ;
  assign n7091 = n7086 & n32629 ;
  assign n7656 = n7087 & n32629 ;
  assign n7657 = n32628 & n7656 ;
  assign n7658 = n7091 | n7657 ;
  assign n7645 = n7641 & n7643 ;
  assign n7646 = n7640 | n7645 ;
  assign n7178 = n6186 & n7162 ;
  assign n7648 = x[126] & n7100 ;
  assign n7649 = x[127] & n7647 ;
  assign n7650 = n7648 | n7649 ;
  assign n7651 = n7178 | n7650 ;
  assign n32630 = ~n7651 ;
  assign n7652 = x[20] & n32630 ;
  assign n7653 = n28114 & n7651 ;
  assign n7654 = n7652 | n7653 ;
  assign n32631 = ~n7654 ;
  assign n7659 = n7646 & n32631 ;
  assign n32632 = ~n7646 ;
  assign n7660 = n32632 & n7654 ;
  assign n7662 = n7659 | n7660 ;
  assign n7663 = n7658 & n7662 ;
  assign n7661 = n7658 | n7660 ;
  assign n8182 = n7659 | n7661 ;
  assign n32633 = ~n7663 ;
  assign n8183 = n32633 & n8182 ;
  assign n32634 = ~n8183 ;
  assign n23175 = n8181 & n32634 ;
  assign n32635 = ~n8181 ;
  assign n23176 = n32635 & n8183 ;
  assign n23177 = n23175 | n23176 ;
  assign n23178 = n23174 & n23177 ;
  assign n27771 = n23174 | n23176 ;
  assign n27772 = n23175 | n27771 ;
  assign n32636 = ~n23178 ;
  assign n211 = n32636 & n27772 ;
  assign n8184 = n8181 & n8183 ;
  assign n23179 = n8184 | n23178 ;
  assign n7655 = n7646 & n7654 ;
  assign n7664 = n7655 | n7663 ;
  assign n7090 = n7085 | n7089 ;
  assign n7143 = x[127] & n7100 ;
  assign n7200 = n5360 & n7162 ;
  assign n7226 = n7143 | n7200 ;
  assign n32637 = ~n7226 ;
  assign n7227 = x[20] & n32637 ;
  assign n7228 = n28114 & n7226 ;
  assign n7229 = n7227 | n7228 ;
  assign n7230 = n7090 | n7229 ;
  assign n7231 = n7090 & n7229 ;
  assign n32638 = ~n7231 ;
  assign n7232 = n7230 & n32638 ;
  assign n5395 = n5302 & n5388 ;
  assign n5277 = x[124] & n5240 ;
  assign n6226 = x[125] & n6179 ;
  assign n6282 = n5277 | n6226 ;
  assign n6283 = x[126] & n5238 ;
  assign n6284 = n6282 | n6283 ;
  assign n6285 = n5395 | n6284 ;
  assign n32639 = ~n6285 ;
  assign n6286 = x[23] & n32639 ;
  assign n6287 = n28221 & n6285 ;
  assign n6288 = n6286 | n6287 ;
  assign n6697 = n6690 | n6696 ;
  assign n6698 = n6288 | n6697 ;
  assign n6699 = n6288 & n6697 ;
  assign n32640 = ~n6699 ;
  assign n6700 = n6698 & n32640 ;
  assign n5421 = n452 & n5417 ;
  assign n382 = x[121] & n330 ;
  assign n417 = x[122] & n390 ;
  assign n5879 = n382 | n417 ;
  assign n5880 = x[123] & n322 ;
  assign n5881 = n5879 | n5880 ;
  assign n5882 = n5421 | n5881 ;
  assign n5883 = x[26] | n5882 ;
  assign n5884 = x[26] & n5882 ;
  assign n32641 = ~n5884 ;
  assign n5885 = n5883 & n32641 ;
  assign n6155 = n5892 & n6153 ;
  assign n6161 = n6155 | n6160 ;
  assign n32642 = ~n6161 ;
  assign n6162 = n5885 & n32642 ;
  assign n32643 = ~n5885 ;
  assign n6164 = n32643 & n6161 ;
  assign n6165 = n6162 | n6164 ;
  assign n4525 = x[118] & n4514 ;
  assign n4601 = x[119] & n4572 ;
  assign n4629 = n4525 | n4601 ;
  assign n4630 = x[120] & n4504 ;
  assign n4631 = n4629 | n4630 ;
  assign n4679 = n4632 & n4678 ;
  assign n4692 = n4631 | n4679 ;
  assign n32644 = ~n4692 ;
  assign n4693 = x[29] & n32644 ;
  assign n4694 = n28483 & n4692 ;
  assign n4695 = n4693 | n4694 ;
  assign n4963 = n4717 & n4961 ;
  assign n4969 = n4963 | n4968 ;
  assign n4970 = n4695 | n4969 ;
  assign n4971 = n4695 & n4969 ;
  assign n32645 = ~n4971 ;
  assign n4972 = n4970 & n32645 ;
  assign n692 = x[115] & n663 ;
  assign n737 = x[116] & n720 ;
  assign n791 = n692 | n737 ;
  assign n792 = x[117] & n652 ;
  assign n793 = n791 | n792 ;
  assign n799 = n779 & n797 ;
  assign n800 = n793 | n799 ;
  assign n801 = x[32] | n800 ;
  assign n802 = x[32] & n800 ;
  assign n32646 = ~n802 ;
  assign n803 = n801 & n32646 ;
  assign n3899 = n3630 & n3897 ;
  assign n4105 = n3901 & n4103 ;
  assign n4106 = n3899 | n4105 ;
  assign n32647 = ~n4106 ;
  assign n4107 = n803 & n32647 ;
  assign n32648 = ~n803 ;
  assign n4294 = n32648 & n4106 ;
  assign n4295 = n4107 | n4294 ;
  assign n4109 = n2887 | n3019 ;
  assign n4110 = n3022 & n3212 ;
  assign n32649 = ~n4110 ;
  assign n4111 = n4109 & n32649 ;
  assign n3878 = n3162 & n3876 ;
  assign n3070 = x[106] & n3031 ;
  assign n3131 = x[107] & n3096 ;
  assign n4112 = n3070 | n3131 ;
  assign n4113 = x[108] & n3027 ;
  assign n4114 = n4112 | n4113 ;
  assign n4115 = n3878 | n4114 ;
  assign n32650 = ~n4115 ;
  assign n4116 = x[41] & n32650 ;
  assign n4117 = n29184 & n4115 ;
  assign n4118 = n4116 | n4117 ;
  assign n32651 = ~n2992 ;
  assign n4119 = n2889 & n32651 ;
  assign n4120 = n3016 | n4119 ;
  assign n3417 = n2635 & n3409 ;
  assign n2516 = x[103] & n2492 ;
  assign n2596 = x[104] & n2557 ;
  assign n4121 = n2516 | n2596 ;
  assign n4122 = x[105] & n2488 ;
  assign n4123 = n4121 | n4122 ;
  assign n4124 = n3417 | n4123 ;
  assign n32652 = ~n4124 ;
  assign n4125 = x[44] & n32652 ;
  assign n4126 = n29400 & n4124 ;
  assign n4127 = n4125 | n4126 ;
  assign n32653 = ~n2970 ;
  assign n4128 = n32653 & n2989 ;
  assign n4129 = n2969 | n4128 ;
  assign n2870 = n2321 & n2867 ;
  assign n2231 = x[100] & n2179 ;
  assign n2276 = x[101] & n2244 ;
  assign n4130 = n2231 | n2276 ;
  assign n4131 = x[102] & n2175 ;
  assign n4132 = n4130 | n4131 ;
  assign n4133 = n2870 | n4132 ;
  assign n32654 = ~n4133 ;
  assign n4134 = x[47] & n32654 ;
  assign n4135 = n29621 & n4133 ;
  assign n4136 = n4134 | n4135 ;
  assign n32655 = ~n2956 ;
  assign n4137 = n32655 & n2963 ;
  assign n4138 = n2955 | n4137 ;
  assign n2316 = n2007 & n2313 ;
  assign n1927 = x[97] & n1866 ;
  assign n1966 = x[98] & n1931 ;
  assign n4139 = n1927 | n1966 ;
  assign n4140 = x[99] & n1862 ;
  assign n4141 = n4139 | n4140 ;
  assign n4142 = n2316 | n4141 ;
  assign n32656 = ~n4142 ;
  assign n4143 = x[50] & n32656 ;
  assign n4144 = n29865 & n4142 ;
  assign n4145 = n4143 | n4144 ;
  assign n32657 = ~n2934 ;
  assign n4146 = n32657 & n2937 ;
  assign n32658 = ~n2940 ;
  assign n4147 = n32658 & n2947 ;
  assign n4148 = n4146 | n4147 ;
  assign n32659 = ~n2906 ;
  assign n4149 = n32659 & n2908 ;
  assign n32660 = ~n2911 ;
  assign n4150 = n32660 & n2918 ;
  assign n4151 = n4149 | n4150 ;
  assign n1484 = n1217 & n1482 ;
  assign n1135 = x[88] & n1079 ;
  assign n1182 = x[89] & n1144 ;
  assign n4152 = n1135 | n1182 ;
  assign n4153 = x[90] & n1075 ;
  assign n4154 = n4152 | n4153 ;
  assign n4155 = n1484 | n4154 ;
  assign n32661 = ~n4155 ;
  assign n4156 = x[59] & n32661 ;
  assign n4157 = n30638 & n4155 ;
  assign n4158 = n4156 | n4157 ;
  assign n32662 = ~n2896 ;
  assign n4159 = n32662 & n2903 ;
  assign n4160 = n2895 | n4159 ;
  assign n27752 = x[83] & n27215 ;
  assign n849 = x[84] & n805 ;
  assign n4161 = n27752 | n849 ;
  assign n4162 = n2892 | n4161 ;
  assign n4164 = n2892 & n4161 ;
  assign n32663 = ~n4164 ;
  assign n4165 = n4162 & n32663 ;
  assign n889 = x[87] & n881 ;
  assign n4166 = x[85] & n900 ;
  assign n4167 = x[86] & n949 ;
  assign n4168 = n4166 | n4167 ;
  assign n4169 = n889 | n4168 ;
  assign n4170 = n1006 & n1522 ;
  assign n4171 = n4169 | n4170 ;
  assign n4172 = n30886 & n4171 ;
  assign n32664 = ~n4171 ;
  assign n4173 = x[62] & n32664 ;
  assign n4174 = n4172 | n4173 ;
  assign n4175 = n4165 | n4174 ;
  assign n4176 = n4165 & n4174 ;
  assign n32665 = ~n4176 ;
  assign n4177 = n4175 & n32665 ;
  assign n32666 = ~n4177 ;
  assign n4178 = n4160 & n32666 ;
  assign n32667 = ~n4160 ;
  assign n4179 = n32667 & n4177 ;
  assign n4180 = n4178 | n4179 ;
  assign n4181 = n4158 | n4180 ;
  assign n4182 = n4158 & n4180 ;
  assign n32668 = ~n4182 ;
  assign n4183 = n4181 & n32668 ;
  assign n4184 = n4151 | n4183 ;
  assign n4185 = n4151 & n4183 ;
  assign n32669 = ~n4185 ;
  assign n4186 = n4184 & n32669 ;
  assign n1687 = n1457 & n1685 ;
  assign n1376 = x[91] & n1319 ;
  assign n1431 = x[92] & n1384 ;
  assign n4187 = n1376 | n1431 ;
  assign n4188 = x[93] & n1315 ;
  assign n4189 = n4187 | n4188 ;
  assign n4190 = n1687 | n4189 ;
  assign n32670 = ~n4190 ;
  assign n4191 = x[56] & n32670 ;
  assign n4192 = n30379 & n4190 ;
  assign n4193 = n4191 | n4192 ;
  assign n4194 = n4186 | n4193 ;
  assign n4195 = n4186 & n4193 ;
  assign n32671 = ~n4195 ;
  assign n4196 = n4194 & n32671 ;
  assign n32672 = ~n2924 ;
  assign n4197 = n32672 & n2931 ;
  assign n32673 = ~n2921 ;
  assign n4198 = n2891 & n32673 ;
  assign n4199 = n4197 | n4198 ;
  assign n32674 = ~n4199 ;
  assign n4200 = n4196 & n32674 ;
  assign n32675 = ~n4196 ;
  assign n4201 = n32675 & n4199 ;
  assign n4202 = n4200 | n4201 ;
  assign n2003 = n1690 & n2000 ;
  assign n1580 = x[94] & n1551 ;
  assign n1646 = x[95] & n1616 ;
  assign n4203 = n1580 | n1646 ;
  assign n4204 = x[96] & n1547 ;
  assign n4205 = n4203 | n4204 ;
  assign n4206 = n2003 | n4205 ;
  assign n32676 = ~n4206 ;
  assign n4207 = x[53] & n32676 ;
  assign n4208 = n30125 & n4206 ;
  assign n4209 = n4207 | n4208 ;
  assign n4210 = n4202 | n4209 ;
  assign n4211 = n4202 & n4209 ;
  assign n32677 = ~n4211 ;
  assign n4212 = n4210 & n32677 ;
  assign n32678 = ~n4148 ;
  assign n4213 = n32678 & n4212 ;
  assign n32679 = ~n4212 ;
  assign n4214 = n4148 & n32679 ;
  assign n4215 = n4213 | n4214 ;
  assign n4216 = n4145 | n4215 ;
  assign n4217 = n4145 & n4215 ;
  assign n32680 = ~n4217 ;
  assign n4218 = n4216 & n32680 ;
  assign n4219 = n4138 | n4218 ;
  assign n4220 = n4138 & n4218 ;
  assign n32681 = ~n4220 ;
  assign n4221 = n4219 & n32681 ;
  assign n4222 = n4136 | n4221 ;
  assign n4223 = n4136 & n4221 ;
  assign n32682 = ~n4223 ;
  assign n4224 = n4222 & n32682 ;
  assign n4225 = n4129 | n4224 ;
  assign n4226 = n4129 & n4224 ;
  assign n32683 = ~n4226 ;
  assign n4227 = n4225 & n32683 ;
  assign n4228 = n4127 | n4227 ;
  assign n4229 = n4127 & n4227 ;
  assign n32684 = ~n4229 ;
  assign n4230 = n4228 & n32684 ;
  assign n4231 = n4120 | n4230 ;
  assign n4232 = n4120 & n4230 ;
  assign n32685 = ~n4232 ;
  assign n4233 = n4231 & n32685 ;
  assign n4234 = n4118 | n4233 ;
  assign n4235 = n4118 & n4233 ;
  assign n32686 = ~n4235 ;
  assign n4236 = n4234 & n32686 ;
  assign n32687 = ~n4236 ;
  assign n4237 = n4111 & n32687 ;
  assign n32688 = ~n4111 ;
  assign n4238 = n32688 & n4236 ;
  assign n4239 = n4237 | n4238 ;
  assign n3454 = x[109] & n3443 ;
  assign n3544 = x[110] & n3508 ;
  assign n4240 = n3454 | n3544 ;
  assign n4241 = x[111] & n3439 ;
  assign n4242 = n4240 | n4241 ;
  assign n4251 = n3574 & n4246 ;
  assign n4257 = n4242 | n4251 ;
  assign n32689 = ~n4257 ;
  assign n4258 = x[38] & n32689 ;
  assign n4259 = n28996 & n4257 ;
  assign n4260 = n4258 | n4259 ;
  assign n32690 = ~n4260 ;
  assign n4261 = n4239 & n32690 ;
  assign n32691 = ~n4239 ;
  assign n4262 = n32691 & n4260 ;
  assign n4263 = n4261 | n4262 ;
  assign n4264 = n3215 & n3431 ;
  assign n4265 = n3434 & n3627 ;
  assign n4266 = n4264 | n4265 ;
  assign n4267 = n4263 | n4266 ;
  assign n4268 = n4263 & n4266 ;
  assign n32692 = ~n4268 ;
  assign n4269 = n4267 & n32692 ;
  assign n3943 = x[112] & n3910 ;
  assign n4019 = x[113] & n3975 ;
  assign n4270 = n3943 | n4019 ;
  assign n4271 = x[114] & n3906 ;
  assign n4272 = n4270 | n4271 ;
  assign n4282 = n4041 & n4276 ;
  assign n4288 = n4272 | n4282 ;
  assign n32693 = ~n4288 ;
  assign n4289 = x[35] & n32693 ;
  assign n4290 = n28822 & n4288 ;
  assign n4291 = n4289 | n4290 ;
  assign n4293 = n4269 & n4291 ;
  assign n4292 = n4269 | n4291 ;
  assign n4296 = n4292 & n4295 ;
  assign n32694 = ~n4293 ;
  assign n4297 = n32694 & n4296 ;
  assign n32695 = ~n4297 ;
  assign n4298 = n4295 & n32695 ;
  assign n4973 = n4292 & n32695 ;
  assign n4974 = n32694 & n4973 ;
  assign n4975 = n4298 | n4974 ;
  assign n4976 = n4972 | n4975 ;
  assign n4977 = n4972 & n4975 ;
  assign n32696 = ~n4977 ;
  assign n6166 = n4976 & n32696 ;
  assign n32697 = ~n6166 ;
  assign n6167 = n6165 & n32697 ;
  assign n32698 = ~n6165 ;
  assign n6701 = n32698 & n6166 ;
  assign n6702 = n6167 | n6701 ;
  assign n6703 = n6700 | n6702 ;
  assign n6704 = n6700 & n6702 ;
  assign n32699 = ~n6704 ;
  assign n7233 = n6703 & n32699 ;
  assign n32700 = ~n7233 ;
  assign n7234 = n7232 & n32700 ;
  assign n32701 = ~n7232 ;
  assign n7665 = n32701 & n7233 ;
  assign n7666 = n7234 | n7665 ;
  assign n32702 = ~n7664 ;
  assign n7667 = n32702 & n7666 ;
  assign n32703 = ~n7666 ;
  assign n23180 = n7664 & n32703 ;
  assign n23181 = n7667 | n23180 ;
  assign n23182 = n23179 | n23181 ;
  assign n23183 = n23179 & n23181 ;
  assign n32704 = ~n23183 ;
  assign n212 = n23182 & n32704 ;
  assign n6705 = n6699 | n6704 ;
  assign n5639 = n5302 & n5629 ;
  assign n5276 = x[125] & n5240 ;
  assign n6278 = x[126] & n6179 ;
  assign n6706 = n5276 | n6278 ;
  assign n6707 = x[127] & n5238 ;
  assign n6708 = n6706 | n6707 ;
  assign n6709 = n5639 | n6708 ;
  assign n32705 = ~n6709 ;
  assign n6710 = x[23] & n32705 ;
  assign n6711 = n28221 & n6709 ;
  assign n6712 = n6710 | n6711 ;
  assign n32706 = ~n6712 ;
  assign n6713 = n6705 & n32706 ;
  assign n32707 = ~n6705 ;
  assign n6715 = n32707 & n6712 ;
  assign n6716 = n6713 | n6715 ;
  assign n5849 = n452 & n5838 ;
  assign n367 = x[122] & n330 ;
  assign n416 = x[123] & n390 ;
  assign n5872 = n367 | n416 ;
  assign n5873 = x[124] & n322 ;
  assign n5874 = n5872 | n5873 ;
  assign n5875 = n5849 | n5874 ;
  assign n32708 = ~n5875 ;
  assign n5876 = x[26] & n32708 ;
  assign n5877 = n28342 & n5875 ;
  assign n5878 = n5876 | n5877 ;
  assign n6163 = n5885 & n6161 ;
  assign n6168 = n6165 & n6166 ;
  assign n6169 = n6163 | n6168 ;
  assign n6170 = n5878 | n6169 ;
  assign n6171 = n5878 & n6169 ;
  assign n32709 = ~n6171 ;
  assign n6172 = n6170 & n32709 ;
  assign n4978 = n4971 | n4977 ;
  assign n4540 = x[119] & n4514 ;
  assign n4590 = x[120] & n4572 ;
  assign n4979 = n4540 | n4590 ;
  assign n4980 = x[121] & n4504 ;
  assign n4981 = n4979 | n4980 ;
  assign n4992 = n4632 & n4985 ;
  assign n4999 = n4981 | n4992 ;
  assign n32710 = ~n4999 ;
  assign n5000 = x[29] & n32710 ;
  assign n5001 = n28483 & n4999 ;
  assign n5002 = n5000 | n5001 ;
  assign n32711 = ~n5002 ;
  assign n5003 = n4978 & n32711 ;
  assign n32712 = ~n4978 ;
  assign n5004 = n32712 & n5002 ;
  assign n5005 = n5003 | n5004 ;
  assign n687 = x[116] & n663 ;
  assign n734 = x[117] & n720 ;
  assign n776 = n687 | n734 ;
  assign n777 = x[118] & n652 ;
  assign n778 = n776 | n777 ;
  assign n786 = n779 & n784 ;
  assign n787 = n778 | n786 ;
  assign n32713 = ~n787 ;
  assign n788 = x[32] & n32713 ;
  assign n789 = n28658 & n787 ;
  assign n790 = n788 | n789 ;
  assign n4108 = n803 & n4106 ;
  assign n4299 = n4108 | n4297 ;
  assign n4300 = n790 | n4299 ;
  assign n4301 = n790 & n4299 ;
  assign n32714 = ~n4301 ;
  assign n4302 = n4300 & n32714 ;
  assign n4303 = n4268 | n4293 ;
  assign n32715 = ~n4215 ;
  assign n4304 = n4145 & n32715 ;
  assign n4305 = n4214 | n4304 ;
  assign n27757 = x[84] & n27215 ;
  assign n819 = x[85] & n805 ;
  assign n4306 = n27757 | n819 ;
  assign n32716 = ~n4306 ;
  assign n4307 = x[20] & n32716 ;
  assign n4308 = n28114 & n4306 ;
  assign n4309 = n4307 | n4308 ;
  assign n4310 = n4161 | n4309 ;
  assign n4312 = n4161 & n4309 ;
  assign n32717 = ~n4312 ;
  assign n4313 = n4310 & n32717 ;
  assign n1723 = n1006 & n1720 ;
  assign n915 = x[86] & n900 ;
  assign n970 = x[87] & n949 ;
  assign n4314 = n915 | n970 ;
  assign n4315 = x[88] & n881 ;
  assign n4316 = n4314 | n4315 ;
  assign n4317 = n1723 | n4316 ;
  assign n32718 = ~n4317 ;
  assign n4318 = x[62] & n32718 ;
  assign n4319 = n30886 & n4317 ;
  assign n4320 = n4318 | n4319 ;
  assign n32719 = ~n4320 ;
  assign n4321 = n4313 & n32719 ;
  assign n32720 = ~n4313 ;
  assign n4322 = n32720 & n4320 ;
  assign n4323 = n4321 | n4322 ;
  assign n32721 = ~n4161 ;
  assign n4163 = n2892 & n32721 ;
  assign n32722 = ~n4165 ;
  assign n4324 = n32722 & n4174 ;
  assign n4325 = n4163 | n4324 ;
  assign n32723 = ~n4325 ;
  assign n4326 = n4323 & n32723 ;
  assign n32724 = ~n4323 ;
  assign n4327 = n32724 & n4325 ;
  assign n4328 = n4326 | n4327 ;
  assign n2049 = n1217 & n2046 ;
  assign n1129 = x[89] & n1079 ;
  assign n1195 = x[90] & n1144 ;
  assign n4329 = n1129 | n1195 ;
  assign n4330 = x[91] & n1075 ;
  assign n4331 = n4329 | n4330 ;
  assign n4332 = n2049 | n4331 ;
  assign n32725 = ~n4332 ;
  assign n4333 = x[59] & n32725 ;
  assign n4334 = n30638 & n4332 ;
  assign n4335 = n4333 | n4334 ;
  assign n32726 = ~n4335 ;
  assign n4336 = n4328 & n32726 ;
  assign n32727 = ~n4328 ;
  assign n4337 = n32727 & n4335 ;
  assign n4338 = n4336 | n4337 ;
  assign n32728 = ~n4180 ;
  assign n4339 = n4158 & n32728 ;
  assign n4340 = n4178 | n4339 ;
  assign n32729 = ~n4340 ;
  assign n4341 = n4338 & n32729 ;
  assign n32730 = ~n4338 ;
  assign n4342 = n32730 & n4340 ;
  assign n4343 = n4341 | n4342 ;
  assign n2416 = n1457 & n2410 ;
  assign n1366 = x[92] & n1319 ;
  assign n1421 = x[93] & n1384 ;
  assign n4344 = n1366 | n1421 ;
  assign n4345 = x[94] & n1315 ;
  assign n4346 = n4344 | n4345 ;
  assign n4347 = n2416 | n4346 ;
  assign n32731 = ~n4347 ;
  assign n4348 = x[56] & n32731 ;
  assign n4349 = n30379 & n4347 ;
  assign n4350 = n4348 | n4349 ;
  assign n4351 = n4343 | n4350 ;
  assign n4352 = n4343 & n4350 ;
  assign n32732 = ~n4352 ;
  assign n4353 = n4351 & n32732 ;
  assign n32733 = ~n4183 ;
  assign n4354 = n4151 & n32733 ;
  assign n32734 = ~n4186 ;
  assign n4355 = n32734 & n4193 ;
  assign n4356 = n4354 | n4355 ;
  assign n4357 = n4353 | n4356 ;
  assign n4358 = n4353 & n4356 ;
  assign n32735 = ~n4358 ;
  assign n4359 = n4357 & n32735 ;
  assign n2443 = n1690 & n2438 ;
  assign n1566 = x[95] & n1551 ;
  assign n1659 = x[96] & n1616 ;
  assign n4360 = n1566 | n1659 ;
  assign n4361 = x[97] & n1547 ;
  assign n4362 = n4360 | n4361 ;
  assign n4363 = n2443 | n4362 ;
  assign n32736 = ~n4363 ;
  assign n4364 = x[53] & n32736 ;
  assign n4365 = n30125 & n4363 ;
  assign n4366 = n4364 | n4365 ;
  assign n32737 = ~n4202 ;
  assign n4367 = n32737 & n4209 ;
  assign n4368 = n4201 | n4367 ;
  assign n4369 = n4366 | n4368 ;
  assign n4370 = n4366 & n4368 ;
  assign n32738 = ~n4370 ;
  assign n4371 = n4369 & n32738 ;
  assign n32739 = ~n4359 ;
  assign n4372 = n32739 & n4371 ;
  assign n32740 = ~n4371 ;
  assign n4373 = n4359 & n32740 ;
  assign n4374 = n4372 | n4373 ;
  assign n2468 = n2007 & n2466 ;
  assign n1911 = x[98] & n1866 ;
  assign n1967 = x[99] & n1931 ;
  assign n4375 = n1911 | n1967 ;
  assign n4376 = x[100] & n1862 ;
  assign n4377 = n4375 | n4376 ;
  assign n4378 = n2468 | n4377 ;
  assign n32741 = ~n4378 ;
  assign n4379 = x[50] & n32741 ;
  assign n4380 = n29865 & n4378 ;
  assign n4381 = n4379 | n4380 ;
  assign n32742 = ~n4381 ;
  assign n4382 = n4374 & n32742 ;
  assign n32743 = ~n4374 ;
  assign n4383 = n32743 & n4381 ;
  assign n4384 = n4382 | n4383 ;
  assign n4385 = n4305 | n4384 ;
  assign n4386 = n4305 & n4384 ;
  assign n32744 = ~n4386 ;
  assign n4387 = n4385 & n32744 ;
  assign n2628 = n2321 & n2626 ;
  assign n2229 = x[101] & n2179 ;
  assign n2274 = x[102] & n2244 ;
  assign n4388 = n2229 | n2274 ;
  assign n4389 = x[103] & n2175 ;
  assign n4390 = n4388 | n4389 ;
  assign n4391 = n2628 | n4390 ;
  assign n32745 = ~n4391 ;
  assign n4392 = x[47] & n32745 ;
  assign n4393 = n29621 & n4391 ;
  assign n4394 = n4392 | n4393 ;
  assign n4395 = n4387 | n4394 ;
  assign n4396 = n4387 & n4394 ;
  assign n32746 = ~n4396 ;
  assign n4397 = n4395 & n32746 ;
  assign n32747 = ~n4218 ;
  assign n4398 = n4138 & n32747 ;
  assign n32748 = ~n4221 ;
  assign n4399 = n4136 & n32748 ;
  assign n4400 = n4398 | n4399 ;
  assign n32749 = ~n4400 ;
  assign n4401 = n4397 & n32749 ;
  assign n32750 = ~n4397 ;
  assign n4402 = n32750 & n4400 ;
  assign n4403 = n4401 | n4402 ;
  assign n3228 = n2635 & n3223 ;
  assign n2515 = x[104] & n2492 ;
  assign n2595 = x[105] & n2557 ;
  assign n4404 = n2515 | n2595 ;
  assign n4405 = x[106] & n2488 ;
  assign n4406 = n4404 | n4405 ;
  assign n4407 = n3228 | n4406 ;
  assign n32751 = ~n4407 ;
  assign n4408 = x[44] & n32751 ;
  assign n4409 = n29400 & n4407 ;
  assign n4410 = n4408 | n4409 ;
  assign n4411 = n4403 | n4410 ;
  assign n4412 = n4403 & n4410 ;
  assign n32752 = ~n4412 ;
  assign n4413 = n4411 & n32752 ;
  assign n32753 = ~n4224 ;
  assign n4414 = n4129 & n32753 ;
  assign n32754 = ~n4227 ;
  assign n4415 = n4127 & n32754 ;
  assign n4416 = n4414 | n4415 ;
  assign n4417 = n4413 | n4416 ;
  assign n4418 = n4413 & n4416 ;
  assign n32755 = ~n4418 ;
  assign n4419 = n4417 & n32755 ;
  assign n3646 = n3162 & n3639 ;
  assign n3057 = x[107] & n3031 ;
  assign n3129 = x[108] & n3096 ;
  assign n4420 = n3057 | n3129 ;
  assign n4421 = x[109] & n3027 ;
  assign n4422 = n4420 | n4421 ;
  assign n4423 = n3646 | n4422 ;
  assign n32756 = ~n4423 ;
  assign n4424 = x[41] & n32756 ;
  assign n4425 = n29184 & n4423 ;
  assign n4426 = n4424 | n4425 ;
  assign n4427 = n4419 | n4426 ;
  assign n4428 = n4419 & n4426 ;
  assign n32757 = ~n4428 ;
  assign n4429 = n4427 & n32757 ;
  assign n32758 = ~n4230 ;
  assign n4430 = n4120 & n32758 ;
  assign n32759 = ~n4233 ;
  assign n4431 = n4118 & n32759 ;
  assign n4432 = n4430 | n4431 ;
  assign n4433 = n4429 | n4432 ;
  assign n4434 = n4429 & n4432 ;
  assign n32760 = ~n4434 ;
  assign n4435 = n4433 & n32760 ;
  assign n3460 = x[110] & n3443 ;
  assign n3532 = x[111] & n3508 ;
  assign n4436 = n3460 | n3532 ;
  assign n4437 = x[112] & n3439 ;
  assign n4438 = n4436 | n4437 ;
  assign n4447 = n3574 & n4442 ;
  assign n4455 = n4438 | n4447 ;
  assign n32761 = ~n4455 ;
  assign n4456 = x[38] & n32761 ;
  assign n4457 = n28996 & n4455 ;
  assign n4458 = n4456 | n4457 ;
  assign n4459 = n4435 | n4458 ;
  assign n4460 = n4435 & n4458 ;
  assign n32762 = ~n4460 ;
  assign n4461 = n4459 & n32762 ;
  assign n4462 = n4111 | n4236 ;
  assign n4463 = n4239 & n4260 ;
  assign n32763 = ~n4463 ;
  assign n4464 = n4462 & n32763 ;
  assign n32764 = ~n4461 ;
  assign n4465 = n32764 & n4464 ;
  assign n32765 = ~n4464 ;
  assign n4466 = n4461 & n32765 ;
  assign n4467 = n4465 | n4466 ;
  assign n3968 = x[113] & n3910 ;
  assign n4017 = x[114] & n3975 ;
  assign n4468 = n3968 | n4017 ;
  assign n4469 = x[115] & n3906 ;
  assign n4470 = n4468 | n4469 ;
  assign n4475 = n4041 & n4474 ;
  assign n4487 = n4470 | n4475 ;
  assign n32766 = ~n4487 ;
  assign n4488 = x[35] & n32766 ;
  assign n4489 = n28822 & n4487 ;
  assign n4490 = n4488 | n4489 ;
  assign n4492 = n4467 & n4490 ;
  assign n4491 = n4467 | n4490 ;
  assign n4493 = n4303 & n4491 ;
  assign n32767 = ~n4492 ;
  assign n4494 = n32767 & n4493 ;
  assign n32768 = ~n4494 ;
  assign n4496 = n4303 & n32768 ;
  assign n4495 = n4492 | n4493 ;
  assign n32769 = ~n4495 ;
  assign n4497 = n4491 & n32769 ;
  assign n4498 = n4496 | n4497 ;
  assign n4499 = n4302 & n4498 ;
  assign n5006 = n4302 | n4498 ;
  assign n5007 = n5005 & n5006 ;
  assign n32770 = ~n4499 ;
  assign n5008 = n32770 & n5007 ;
  assign n32771 = ~n5008 ;
  assign n6173 = n5005 & n32771 ;
  assign n6174 = n5006 & n32771 ;
  assign n6175 = n32770 & n6174 ;
  assign n6176 = n6173 | n6175 ;
  assign n6177 = n6172 & n6176 ;
  assign n6717 = n6172 | n6176 ;
  assign n6718 = n6716 & n6717 ;
  assign n32772 = ~n6177 ;
  assign n6719 = n32772 & n6718 ;
  assign n32773 = ~n6719 ;
  assign n6725 = n6716 & n32773 ;
  assign n6726 = n6717 & n32773 ;
  assign n6727 = n32772 & n6726 ;
  assign n6728 = n6725 | n6727 ;
  assign n7235 = n7232 & n7233 ;
  assign n7236 = n7231 | n7235 ;
  assign n7237 = n6728 | n7236 ;
  assign n7238 = n6728 & n7236 ;
  assign n32774 = ~n7238 ;
  assign n7239 = n7237 & n32774 ;
  assign n7668 = n7664 & n7666 ;
  assign n23184 = n7668 | n23183 ;
  assign n23185 = n7239 & n23184 ;
  assign n27775 = n7239 | n23184 ;
  assign n32775 = ~n23185 ;
  assign n213 = n32775 & n27775 ;
  assign n6178 = n6171 | n6177 ;
  assign n6180 = x[126] & n5240 ;
  assign n6181 = x[127] & n6179 ;
  assign n6182 = n6180 | n6181 ;
  assign n6194 = n5302 & n6186 ;
  assign n6201 = n6182 | n6194 ;
  assign n32776 = ~n6201 ;
  assign n6202 = x[23] & n32776 ;
  assign n6203 = n28221 & n6201 ;
  assign n6204 = n6202 | n6203 ;
  assign n32777 = ~n6204 ;
  assign n6205 = n6178 & n32777 ;
  assign n32778 = ~n6178 ;
  assign n6207 = n32778 & n6204 ;
  assign n6208 = n6205 | n6207 ;
  assign n375 = x[123] & n330 ;
  assign n409 = x[124] & n390 ;
  assign n449 = n375 | n409 ;
  assign n450 = x[125] & n322 ;
  assign n451 = n449 | n450 ;
  assign n643 = n452 & n642 ;
  assign n644 = n451 | n643 ;
  assign n32779 = ~n644 ;
  assign n645 = x[26] & n32779 ;
  assign n646 = n28342 & n644 ;
  assign n647 = n645 | n646 ;
  assign n5009 = n4978 & n5002 ;
  assign n5010 = n5008 | n5009 ;
  assign n5011 = n647 | n5010 ;
  assign n5012 = n647 & n5010 ;
  assign n32780 = ~n5012 ;
  assign n5013 = n5011 & n32780 ;
  assign n5014 = n4301 | n4499 ;
  assign n4505 = x[122] & n4504 ;
  assign n5015 = x[120] & n4514 ;
  assign n5016 = x[121] & n4572 ;
  assign n5017 = n5015 | n5016 ;
  assign n5018 = n4505 | n5017 ;
  assign n5033 = n4632 & n5022 ;
  assign n5034 = n5018 | n5033 ;
  assign n5035 = n28483 & n5034 ;
  assign n32781 = ~n5034 ;
  assign n5036 = x[29] & n32781 ;
  assign n5037 = n5035 | n5036 ;
  assign n5038 = n5014 | n5037 ;
  assign n5039 = n5014 & n5037 ;
  assign n32782 = ~n5039 ;
  assign n5040 = n5038 & n32782 ;
  assign n695 = x[117] & n663 ;
  assign n750 = x[118] & n720 ;
  assign n5041 = n695 | n750 ;
  assign n5042 = x[119] & n652 ;
  assign n5043 = n5041 | n5042 ;
  assign n5055 = n779 & n5047 ;
  assign n5061 = n5043 | n5055 ;
  assign n32783 = ~n5061 ;
  assign n5062 = x[32] & n32783 ;
  assign n5063 = n28658 & n5061 ;
  assign n5064 = n5062 | n5063 ;
  assign n32784 = ~n5064 ;
  assign n5065 = n4495 & n32784 ;
  assign n5066 = n32769 & n5064 ;
  assign n5067 = n5065 | n5066 ;
  assign n32785 = ~n4387 ;
  assign n5068 = n32785 & n4394 ;
  assign n5069 = n4402 | n5068 ;
  assign n3005 = n2321 & n3001 ;
  assign n2216 = x[102] & n2179 ;
  assign n2285 = x[103] & n2244 ;
  assign n5149 = n2216 | n2285 ;
  assign n5150 = x[104] & n2175 ;
  assign n5151 = n5149 | n5150 ;
  assign n5152 = n3005 | n5151 ;
  assign n5153 = x[47] | n5152 ;
  assign n5154 = x[47] & n5152 ;
  assign n32786 = ~n5154 ;
  assign n5155 = n5153 & n32786 ;
  assign n32787 = ~n4384 ;
  assign n5070 = n4305 & n32787 ;
  assign n5071 = n4383 | n5070 ;
  assign n5072 = n4337 | n4342 ;
  assign n1844 = n1217 & n1841 ;
  assign n1110 = x[90] & n1079 ;
  assign n1198 = x[91] & n1144 ;
  assign n5073 = n1110 | n1198 ;
  assign n5074 = x[92] & n1075 ;
  assign n5075 = n5073 | n5074 ;
  assign n5076 = n1844 | n5075 ;
  assign n5077 = x[59] | n5076 ;
  assign n5078 = x[59] & n5076 ;
  assign n32788 = ~n5078 ;
  assign n5079 = n5077 & n32788 ;
  assign n5080 = n4322 | n4327 ;
  assign n27767 = x[85] & n27215 ;
  assign n810 = x[86] & n805 ;
  assign n5081 = n27767 | n810 ;
  assign n32789 = ~n4309 ;
  assign n4311 = n4161 & n32789 ;
  assign n5082 = n4308 | n4311 ;
  assign n5083 = n5081 | n5082 ;
  assign n5084 = n5081 & n5082 ;
  assign n32790 = ~n5084 ;
  assign n5085 = n5083 & n32790 ;
  assign n892 = x[89] & n881 ;
  assign n5086 = x[87] & n900 ;
  assign n5087 = x[88] & n949 ;
  assign n5088 = n5086 | n5087 ;
  assign n5089 = n892 | n5088 ;
  assign n5090 = n1006 & n1453 ;
  assign n5091 = n5089 | n5090 ;
  assign n5092 = n30886 & n5091 ;
  assign n32791 = ~n5091 ;
  assign n5093 = x[62] & n32791 ;
  assign n5094 = n5092 | n5093 ;
  assign n5095 = n5085 | n5094 ;
  assign n5096 = n5085 & n5094 ;
  assign n32792 = ~n5096 ;
  assign n5097 = n5095 & n32792 ;
  assign n32793 = ~n5097 ;
  assign n5098 = n5080 & n32793 ;
  assign n32794 = ~n5080 ;
  assign n5099 = n32794 & n5097 ;
  assign n5100 = n5098 | n5099 ;
  assign n32795 = ~n5100 ;
  assign n5101 = n5079 & n32795 ;
  assign n32796 = ~n5079 ;
  assign n5102 = n32796 & n5100 ;
  assign n5103 = n5101 | n5102 ;
  assign n5104 = n5072 | n5103 ;
  assign n5105 = n5072 & n5103 ;
  assign n32797 = ~n5105 ;
  assign n5106 = n5104 & n32797 ;
  assign n2154 = n1457 & n2152 ;
  assign n1368 = x[93] & n1319 ;
  assign n1434 = x[94] & n1384 ;
  assign n5107 = n1368 | n1434 ;
  assign n5108 = x[95] & n1315 ;
  assign n5109 = n5107 | n5108 ;
  assign n5110 = n2154 | n5109 ;
  assign n32798 = ~n5110 ;
  assign n5111 = x[56] & n32798 ;
  assign n5112 = n30379 & n5110 ;
  assign n5113 = n5111 | n5112 ;
  assign n5114 = n5106 | n5113 ;
  assign n5115 = n5106 & n5113 ;
  assign n32799 = ~n5115 ;
  assign n5116 = n5114 & n32799 ;
  assign n32800 = ~n4343 ;
  assign n5117 = n32800 & n4350 ;
  assign n32801 = ~n4353 ;
  assign n5118 = n32801 & n4356 ;
  assign n5119 = n5117 | n5118 ;
  assign n32802 = ~n5119 ;
  assign n5120 = n5116 & n32802 ;
  assign n32803 = ~n5116 ;
  assign n5121 = n32803 & n5119 ;
  assign n5122 = n5120 | n5121 ;
  assign n2844 = n1690 & n2841 ;
  assign n1600 = x[96] & n1551 ;
  assign n1669 = x[97] & n1616 ;
  assign n5123 = n1600 | n1669 ;
  assign n5124 = x[98] & n1547 ;
  assign n5125 = n5123 | n5124 ;
  assign n5126 = n2844 | n5125 ;
  assign n32804 = ~n5126 ;
  assign n5127 = x[53] & n32804 ;
  assign n5128 = n30125 & n5126 ;
  assign n5129 = n5127 | n5128 ;
  assign n5130 = n5122 | n5129 ;
  assign n5131 = n5122 & n5129 ;
  assign n32805 = ~n5131 ;
  assign n5132 = n5130 & n32805 ;
  assign n5133 = n4370 | n4372 ;
  assign n5134 = n5132 | n5133 ;
  assign n5135 = n5132 & n5133 ;
  assign n32806 = ~n5135 ;
  assign n5136 = n5134 & n32806 ;
  assign n2978 = n2007 & n2977 ;
  assign n1874 = x[99] & n1866 ;
  assign n1968 = x[100] & n1931 ;
  assign n5137 = n1874 | n1968 ;
  assign n5138 = x[101] & n1862 ;
  assign n5139 = n5137 | n5138 ;
  assign n5140 = n2978 | n5139 ;
  assign n32807 = ~n5140 ;
  assign n5141 = x[50] & n32807 ;
  assign n5142 = n29865 & n5140 ;
  assign n5143 = n5141 | n5142 ;
  assign n5144 = n5136 | n5143 ;
  assign n5145 = n5136 & n5143 ;
  assign n32808 = ~n5145 ;
  assign n5146 = n5144 & n32808 ;
  assign n5147 = n5071 | n5146 ;
  assign n5148 = n5071 & n5146 ;
  assign n32809 = ~n5148 ;
  assign n5156 = n5147 & n32809 ;
  assign n32810 = ~n5156 ;
  assign n5157 = n5155 & n32810 ;
  assign n32811 = ~n5155 ;
  assign n5158 = n5147 & n32811 ;
  assign n5159 = n32809 & n5158 ;
  assign n5160 = n5157 | n5159 ;
  assign n32812 = ~n5069 ;
  assign n5161 = n32812 & n5160 ;
  assign n32813 = ~n5160 ;
  assign n5162 = n5069 & n32813 ;
  assign n5163 = n5161 | n5162 ;
  assign n3202 = n2635 & n3199 ;
  assign n2529 = x[105] & n2492 ;
  assign n2562 = x[106] & n2557 ;
  assign n5164 = n2529 | n2562 ;
  assign n5165 = x[107] & n2488 ;
  assign n5166 = n5164 | n5165 ;
  assign n5167 = n3202 | n5166 ;
  assign n32814 = ~n5167 ;
  assign n5168 = x[44] & n32814 ;
  assign n5169 = n29400 & n5167 ;
  assign n5170 = n5168 | n5169 ;
  assign n5171 = n5163 | n5170 ;
  assign n5172 = n5163 & n5170 ;
  assign n32815 = ~n5172 ;
  assign n5173 = n5171 & n32815 ;
  assign n32816 = ~n4403 ;
  assign n5174 = n32816 & n4410 ;
  assign n32817 = ~n4413 ;
  assign n5175 = n32817 & n4416 ;
  assign n5176 = n5174 | n5175 ;
  assign n5177 = n5173 | n5176 ;
  assign n5178 = n5173 & n5176 ;
  assign n32818 = ~n5178 ;
  assign n5179 = n5177 & n32818 ;
  assign n3619 = n3162 & n3615 ;
  assign n3088 = x[108] & n3031 ;
  assign n3156 = x[109] & n3096 ;
  assign n5180 = n3088 | n3156 ;
  assign n5181 = x[110] & n3027 ;
  assign n5182 = n5180 | n5181 ;
  assign n5183 = n3619 | n5182 ;
  assign n32819 = ~n5183 ;
  assign n5184 = x[41] & n32819 ;
  assign n5185 = n29184 & n5183 ;
  assign n5186 = n5184 | n5185 ;
  assign n5187 = n5179 | n5186 ;
  assign n5188 = n5179 & n5186 ;
  assign n32820 = ~n5188 ;
  assign n5189 = n5187 & n32820 ;
  assign n32821 = ~n4419 ;
  assign n5190 = n32821 & n4426 ;
  assign n32822 = ~n4429 ;
  assign n5191 = n32822 & n4432 ;
  assign n5192 = n5190 | n5191 ;
  assign n32823 = ~n5192 ;
  assign n5193 = n5189 & n32823 ;
  assign n32824 = ~n5189 ;
  assign n5194 = n32824 & n5192 ;
  assign n5195 = n5193 | n5194 ;
  assign n4092 = n3574 & n4087 ;
  assign n3493 = x[111] & n3443 ;
  assign n3530 = x[112] & n3508 ;
  assign n5196 = n3493 | n3530 ;
  assign n5197 = x[113] & n3439 ;
  assign n5198 = n5196 | n5197 ;
  assign n5199 = n4092 | n5198 ;
  assign n32825 = ~n5199 ;
  assign n5200 = x[38] & n32825 ;
  assign n5201 = n28996 & n5199 ;
  assign n5202 = n5200 | n5201 ;
  assign n5203 = n5195 | n5202 ;
  assign n5204 = n5195 & n5202 ;
  assign n32826 = ~n5204 ;
  assign n5205 = n5203 & n32826 ;
  assign n32827 = ~n4435 ;
  assign n5206 = n32827 & n4458 ;
  assign n5207 = n4461 | n4464 ;
  assign n32828 = ~n5206 ;
  assign n5208 = n32828 & n5207 ;
  assign n32829 = ~n5205 ;
  assign n5209 = n32829 & n5208 ;
  assign n32830 = ~n5208 ;
  assign n5210 = n5205 & n32830 ;
  assign n5211 = n5209 | n5210 ;
  assign n4708 = n4041 & n4702 ;
  assign n3939 = x[114] & n3910 ;
  assign n4031 = x[115] & n3975 ;
  assign n5212 = n3939 | n4031 ;
  assign n5213 = x[116] & n3906 ;
  assign n5214 = n5212 | n5213 ;
  assign n5215 = n4708 | n5214 ;
  assign n32831 = ~n5215 ;
  assign n5216 = x[35] & n32831 ;
  assign n5217 = n28822 & n5215 ;
  assign n5218 = n5216 | n5217 ;
  assign n32832 = ~n5218 ;
  assign n5219 = n5211 & n32832 ;
  assign n32833 = ~n5211 ;
  assign n5220 = n32833 & n5218 ;
  assign n5221 = n5219 | n5220 ;
  assign n5222 = n5067 & n5221 ;
  assign n5223 = n5067 | n5221 ;
  assign n5224 = n5040 & n5223 ;
  assign n32834 = ~n5222 ;
  assign n5225 = n32834 & n5224 ;
  assign n32835 = ~n5225 ;
  assign n5226 = n5040 & n32835 ;
  assign n5227 = n5223 & n32835 ;
  assign n5228 = n32834 & n5227 ;
  assign n5229 = n5226 | n5228 ;
  assign n5230 = n5013 & n5229 ;
  assign n6209 = n5013 | n5229 ;
  assign n6210 = n6208 & n6209 ;
  assign n32836 = ~n5230 ;
  assign n6211 = n32836 & n6210 ;
  assign n32837 = ~n6211 ;
  assign n6217 = n6208 & n32837 ;
  assign n6216 = n6209 & n32837 ;
  assign n6218 = n32836 & n6216 ;
  assign n6219 = n6217 | n6218 ;
  assign n6714 = n6705 & n6712 ;
  assign n6720 = n6714 | n6719 ;
  assign n32838 = ~n6720 ;
  assign n6721 = n6219 & n32838 ;
  assign n32839 = ~n6219 ;
  assign n6723 = n32839 & n6720 ;
  assign n6724 = n6721 | n6723 ;
  assign n23186 = n7238 | n23185 ;
  assign n23187 = n6724 | n23186 ;
  assign n23188 = n6724 & n23186 ;
  assign n32840 = ~n23188 ;
  assign n214 = n23187 & n32840 ;
  assign n6722 = n6219 & n6720 ;
  assign n23189 = n6722 | n23188 ;
  assign n6206 = n6178 & n6204 ;
  assign n6212 = n6206 | n6211 ;
  assign n5231 = n5012 | n5230 ;
  assign n5284 = x[127] & n5240 ;
  assign n5367 = n5302 & n5360 ;
  assign n5375 = n5284 | n5367 ;
  assign n32841 = ~n5375 ;
  assign n5376 = x[23] & n32841 ;
  assign n5377 = n28221 & n5375 ;
  assign n5378 = n5376 | n5377 ;
  assign n5379 = n5231 | n5378 ;
  assign n5380 = n5231 & n5378 ;
  assign n32842 = ~n5380 ;
  assign n5381 = n5379 & n32842 ;
  assign n371 = x[124] & n330 ;
  assign n407 = x[125] & n390 ;
  assign n5382 = n371 | n407 ;
  assign n5383 = x[126] & n322 ;
  assign n5384 = n5382 | n5383 ;
  assign n5399 = n452 & n5388 ;
  assign n5403 = n5384 | n5399 ;
  assign n32843 = ~n5403 ;
  assign n5404 = x[26] & n32843 ;
  assign n5405 = n28342 & n5403 ;
  assign n5406 = n5404 | n5405 ;
  assign n5407 = n5039 | n5225 ;
  assign n5408 = n5406 | n5407 ;
  assign n5409 = n5406 & n5407 ;
  assign n32844 = ~n5409 ;
  assign n5410 = n5408 & n32844 ;
  assign n4539 = x[121] & n4514 ;
  assign n4595 = x[122] & n4572 ;
  assign n5411 = n4539 | n4595 ;
  assign n5412 = x[123] & n4504 ;
  assign n5413 = n5411 | n5412 ;
  assign n5424 = n4632 & n5417 ;
  assign n5432 = n5413 | n5424 ;
  assign n32845 = ~n5432 ;
  assign n5433 = x[29] & n32845 ;
  assign n5434 = n28483 & n5432 ;
  assign n5435 = n5433 | n5434 ;
  assign n5436 = n4495 & n5064 ;
  assign n5437 = n5222 | n5436 ;
  assign n5438 = n5435 | n5437 ;
  assign n5439 = n5435 & n5437 ;
  assign n32846 = ~n5439 ;
  assign n5440 = n5438 & n32846 ;
  assign n4684 = n779 & n4678 ;
  assign n688 = x[118] & n663 ;
  assign n747 = x[119] & n720 ;
  assign n5441 = n688 | n747 ;
  assign n5442 = x[120] & n652 ;
  assign n5443 = n5441 | n5442 ;
  assign n5444 = n4684 | n5443 ;
  assign n5445 = x[32] | n5444 ;
  assign n5446 = x[32] & n5444 ;
  assign n32847 = ~n5446 ;
  assign n5447 = n5445 & n32847 ;
  assign n5448 = n5205 | n5208 ;
  assign n5449 = n5211 & n5218 ;
  assign n32848 = ~n5449 ;
  assign n5450 = n5448 & n32848 ;
  assign n5451 = n5447 & n5450 ;
  assign n5452 = n5447 | n5450 ;
  assign n32849 = ~n5451 ;
  assign n5453 = n32849 & n5452 ;
  assign n4061 = n797 & n4041 ;
  assign n3949 = x[115] & n3910 ;
  assign n4009 = x[116] & n3975 ;
  assign n5454 = n3949 | n4009 ;
  assign n5455 = x[117] & n3906 ;
  assign n5456 = n5454 | n5455 ;
  assign n5457 = n4061 | n5456 ;
  assign n5458 = x[35] | n5457 ;
  assign n5459 = x[35] & n5457 ;
  assign n32850 = ~n5459 ;
  assign n5460 = n5458 & n32850 ;
  assign n32851 = ~n5195 ;
  assign n5461 = n32851 & n5202 ;
  assign n5462 = n5194 | n5461 ;
  assign n32852 = ~n5163 ;
  assign n5463 = n32852 & n5170 ;
  assign n5464 = n5162 | n5463 ;
  assign n3877 = n2635 & n3876 ;
  assign n2530 = x[106] & n2492 ;
  assign n2589 = x[107] & n2557 ;
  assign n5465 = n2530 | n2589 ;
  assign n5466 = x[108] & n2488 ;
  assign n5467 = n5465 | n5466 ;
  assign n5468 = n3877 | n5467 ;
  assign n32853 = ~n5468 ;
  assign n5469 = x[44] & n32853 ;
  assign n5470 = n29400 & n5468 ;
  assign n5471 = n5469 | n5470 ;
  assign n32854 = ~n5146 ;
  assign n5472 = n5071 & n32854 ;
  assign n5473 = n5157 | n5472 ;
  assign n32855 = ~n5122 ;
  assign n5474 = n32855 & n5129 ;
  assign n5475 = n5121 | n5474 ;
  assign n2315 = n1690 & n2313 ;
  assign n1601 = x[97] & n1551 ;
  assign n1640 = x[98] & n1616 ;
  assign n5476 = n1601 | n1640 ;
  assign n5477 = x[99] & n1547 ;
  assign n5478 = n5476 | n5477 ;
  assign n5479 = n2315 | n5478 ;
  assign n32856 = ~n5479 ;
  assign n5480 = x[53] & n32856 ;
  assign n5481 = n30125 & n5479 ;
  assign n5482 = n5480 | n5481 ;
  assign n32857 = ~n5103 ;
  assign n5483 = n5072 & n32857 ;
  assign n32858 = ~n5106 ;
  assign n5484 = n32858 & n5113 ;
  assign n5485 = n5483 | n5484 ;
  assign n32859 = ~n5081 ;
  assign n5486 = n32859 & n5082 ;
  assign n32860 = ~n5085 ;
  assign n5487 = n32860 & n5094 ;
  assign n5488 = n5486 | n5487 ;
  assign n27776 = x[86] & n27215 ;
  assign n855 = x[87] & n805 ;
  assign n5489 = n27776 | n855 ;
  assign n5490 = n5081 | n5489 ;
  assign n5491 = n5081 & n5489 ;
  assign n32861 = ~n5491 ;
  assign n5492 = n5490 & n32861 ;
  assign n887 = x[90] & n881 ;
  assign n5493 = x[88] & n900 ;
  assign n5494 = x[89] & n949 ;
  assign n5495 = n5493 | n5494 ;
  assign n5496 = n887 | n5495 ;
  assign n5497 = n1006 & n1482 ;
  assign n5498 = n5496 | n5497 ;
  assign n5499 = n30886 & n5498 ;
  assign n32862 = ~n5498 ;
  assign n5500 = x[62] & n32862 ;
  assign n5501 = n5499 | n5500 ;
  assign n5502 = n5492 | n5501 ;
  assign n5503 = n5492 & n5501 ;
  assign n32863 = ~n5503 ;
  assign n5504 = n5502 & n32863 ;
  assign n5505 = n5488 | n5504 ;
  assign n5506 = n5488 & n5504 ;
  assign n32864 = ~n5506 ;
  assign n5507 = n5505 & n32864 ;
  assign n1689 = n1217 & n1685 ;
  assign n1105 = x[91] & n1079 ;
  assign n1194 = x[92] & n1144 ;
  assign n5508 = n1105 | n1194 ;
  assign n5509 = x[93] & n1075 ;
  assign n5510 = n5508 | n5509 ;
  assign n5511 = n1689 | n5510 ;
  assign n32865 = ~n5511 ;
  assign n5512 = x[59] & n32865 ;
  assign n5513 = n30638 & n5511 ;
  assign n5514 = n5512 | n5513 ;
  assign n5515 = n5507 | n5514 ;
  assign n5516 = n5507 & n5514 ;
  assign n32866 = ~n5516 ;
  assign n5517 = n5515 & n32866 ;
  assign n5518 = n5098 | n5101 ;
  assign n5519 = n5517 | n5518 ;
  assign n5520 = n5517 & n5518 ;
  assign n32867 = ~n5520 ;
  assign n5521 = n5519 & n32867 ;
  assign n2005 = n1457 & n2000 ;
  assign n1330 = x[94] & n1319 ;
  assign n1418 = x[95] & n1384 ;
  assign n5522 = n1330 | n1418 ;
  assign n5523 = x[96] & n1315 ;
  assign n5524 = n5522 | n5523 ;
  assign n5525 = n2005 | n5524 ;
  assign n32868 = ~n5525 ;
  assign n5526 = x[56] & n32868 ;
  assign n5527 = n30379 & n5525 ;
  assign n5528 = n5526 | n5527 ;
  assign n5529 = n5521 | n5528 ;
  assign n5530 = n5521 & n5528 ;
  assign n32869 = ~n5530 ;
  assign n5531 = n5529 & n32869 ;
  assign n5532 = n5485 | n5531 ;
  assign n5533 = n5485 & n5531 ;
  assign n32870 = ~n5533 ;
  assign n5534 = n5532 & n32870 ;
  assign n5535 = n5482 | n5534 ;
  assign n5536 = n5482 & n5534 ;
  assign n32871 = ~n5536 ;
  assign n5537 = n5535 & n32871 ;
  assign n5538 = n5475 | n5537 ;
  assign n5539 = n5475 & n5537 ;
  assign n32872 = ~n5539 ;
  assign n5540 = n5538 & n32872 ;
  assign n2872 = n2007 & n2867 ;
  assign n1912 = x[100] & n1866 ;
  assign n1978 = x[101] & n1931 ;
  assign n5541 = n1912 | n1978 ;
  assign n5542 = x[102] & n1862 ;
  assign n5543 = n5541 | n5542 ;
  assign n5544 = n2872 | n5543 ;
  assign n32873 = ~n5544 ;
  assign n5545 = x[50] & n32873 ;
  assign n5546 = n29865 & n5544 ;
  assign n5547 = n5545 | n5546 ;
  assign n5548 = n5540 | n5547 ;
  assign n5549 = n5540 & n5547 ;
  assign n32874 = ~n5549 ;
  assign n5550 = n5548 & n32874 ;
  assign n32875 = ~n5132 ;
  assign n5551 = n32875 & n5133 ;
  assign n32876 = ~n5136 ;
  assign n5552 = n32876 & n5143 ;
  assign n5553 = n5551 | n5552 ;
  assign n32877 = ~n5553 ;
  assign n5554 = n5550 & n32877 ;
  assign n32878 = ~n5550 ;
  assign n5555 = n32878 & n5553 ;
  assign n5556 = n5554 | n5555 ;
  assign n3416 = n2321 & n3409 ;
  assign n2197 = x[103] & n2179 ;
  assign n2253 = x[104] & n2244 ;
  assign n5557 = n2197 | n2253 ;
  assign n5558 = x[105] & n2175 ;
  assign n5559 = n5557 | n5558 ;
  assign n5560 = n3416 | n5559 ;
  assign n32879 = ~n5560 ;
  assign n5561 = x[47] & n32879 ;
  assign n5562 = n29621 & n5560 ;
  assign n5563 = n5561 | n5562 ;
  assign n32880 = ~n5563 ;
  assign n5564 = n5556 & n32880 ;
  assign n32881 = ~n5556 ;
  assign n5565 = n32881 & n5563 ;
  assign n5566 = n5564 | n5565 ;
  assign n32882 = ~n5473 ;
  assign n5567 = n32882 & n5566 ;
  assign n32883 = ~n5566 ;
  assign n5568 = n5473 & n32883 ;
  assign n5569 = n5567 | n5568 ;
  assign n5570 = n5471 | n5569 ;
  assign n5571 = n5471 & n5569 ;
  assign n32884 = ~n5571 ;
  assign n5572 = n5570 & n32884 ;
  assign n5573 = n5464 | n5572 ;
  assign n5574 = n5464 & n5572 ;
  assign n32885 = ~n5574 ;
  assign n5575 = n5573 & n32885 ;
  assign n4249 = n3162 & n4246 ;
  assign n3072 = x[109] & n3031 ;
  assign n3140 = x[110] & n3096 ;
  assign n5576 = n3072 | n3140 ;
  assign n5577 = x[111] & n3027 ;
  assign n5578 = n5576 | n5577 ;
  assign n5579 = n4249 | n5578 ;
  assign n32886 = ~n5579 ;
  assign n5580 = x[41] & n32886 ;
  assign n5581 = n29184 & n5579 ;
  assign n5582 = n5580 | n5581 ;
  assign n5583 = n5575 | n5582 ;
  assign n5584 = n5575 & n5582 ;
  assign n32887 = ~n5584 ;
  assign n5585 = n5583 & n32887 ;
  assign n32888 = ~n5173 ;
  assign n5586 = n32888 & n5176 ;
  assign n32889 = ~n5179 ;
  assign n5587 = n32889 & n5186 ;
  assign n5588 = n5586 | n5587 ;
  assign n32890 = ~n5588 ;
  assign n5589 = n5585 & n32890 ;
  assign n32891 = ~n5585 ;
  assign n5590 = n32891 & n5588 ;
  assign n5591 = n5589 | n5590 ;
  assign n4279 = n3574 & n4276 ;
  assign n3484 = x[112] & n3443 ;
  assign n3549 = x[113] & n3508 ;
  assign n5592 = n3484 | n3549 ;
  assign n5593 = x[114] & n3439 ;
  assign n5594 = n5592 | n5593 ;
  assign n5595 = n4279 | n5594 ;
  assign n32892 = ~n5595 ;
  assign n5596 = x[38] & n32892 ;
  assign n5597 = n28996 & n5595 ;
  assign n5598 = n5596 | n5597 ;
  assign n5599 = n5591 | n5598 ;
  assign n5600 = n5591 & n5598 ;
  assign n32893 = ~n5600 ;
  assign n5601 = n5599 & n32893 ;
  assign n5602 = n5462 | n5601 ;
  assign n5603 = n5462 & n5601 ;
  assign n32894 = ~n5603 ;
  assign n5604 = n5602 & n32894 ;
  assign n5605 = n5460 & n5604 ;
  assign n5606 = n5460 | n5604 ;
  assign n32895 = ~n5605 ;
  assign n5607 = n32895 & n5606 ;
  assign n32896 = ~n5453 ;
  assign n5608 = n32896 & n5607 ;
  assign n32897 = ~n5607 ;
  assign n5609 = n5453 & n32897 ;
  assign n5610 = n5608 | n5609 ;
  assign n32898 = ~n5440 ;
  assign n5611 = n32898 & n5610 ;
  assign n32899 = ~n5610 ;
  assign n5612 = n5440 & n32899 ;
  assign n5613 = n5611 | n5612 ;
  assign n32900 = ~n5613 ;
  assign n5614 = n5410 & n32900 ;
  assign n32901 = ~n5410 ;
  assign n5615 = n32901 & n5613 ;
  assign n5616 = n5614 | n5615 ;
  assign n32902 = ~n5616 ;
  assign n5618 = n5381 & n32902 ;
  assign n32903 = ~n5381 ;
  assign n6213 = n32903 & n5616 ;
  assign n6214 = n5618 | n6213 ;
  assign n32904 = ~n6214 ;
  assign n23190 = n6212 & n32904 ;
  assign n32905 = ~n6212 ;
  assign n23191 = n32905 & n6214 ;
  assign n23192 = n23190 | n23191 ;
  assign n23193 = n23189 & n23192 ;
  assign n27778 = n23189 | n23191 ;
  assign n27779 = n23190 | n27778 ;
  assign n32906 = ~n23193 ;
  assign n215 = n32906 & n27779 ;
  assign n6215 = n6212 & n6214 ;
  assign n23194 = n6215 | n23193 ;
  assign n5617 = n5381 & n5616 ;
  assign n5619 = n5380 | n5617 ;
  assign n5620 = n5410 & n5613 ;
  assign n5621 = n5409 | n5620 ;
  assign n363 = x[125] & n330 ;
  assign n427 = x[126] & n390 ;
  assign n5622 = n363 | n427 ;
  assign n5623 = x[127] & n322 ;
  assign n5624 = n5622 | n5623 ;
  assign n5641 = n452 & n5629 ;
  assign n5644 = n5624 | n5641 ;
  assign n32907 = ~n5644 ;
  assign n5645 = x[26] & n32907 ;
  assign n5646 = n28342 & n5644 ;
  assign n5647 = n5645 | n5646 ;
  assign n5648 = n5621 | n5647 ;
  assign n5649 = n5621 & n5647 ;
  assign n32908 = ~n5649 ;
  assign n5650 = n5648 & n32908 ;
  assign n5830 = n5440 & n5610 ;
  assign n5831 = n5439 | n5830 ;
  assign n4524 = x[122] & n4514 ;
  assign n4588 = x[123] & n4572 ;
  assign n5832 = n4524 | n4588 ;
  assign n5833 = x[124] & n4504 ;
  assign n5834 = n5832 | n5833 ;
  assign n5846 = n4632 & n5838 ;
  assign n5853 = n5834 | n5846 ;
  assign n32909 = ~n5853 ;
  assign n5854 = x[29] & n32909 ;
  assign n5855 = n28483 & n5853 ;
  assign n5856 = n5854 | n5855 ;
  assign n5857 = n5831 | n5856 ;
  assign n5858 = n5831 & n5856 ;
  assign n32910 = ~n5858 ;
  assign n5859 = n5857 & n32910 ;
  assign n4987 = n779 & n4985 ;
  assign n697 = x[119] & n663 ;
  assign n743 = x[120] & n720 ;
  assign n5651 = n697 | n743 ;
  assign n5652 = x[121] & n652 ;
  assign n5653 = n5651 | n5652 ;
  assign n5654 = n4987 | n5653 ;
  assign n5655 = x[32] | n5654 ;
  assign n5656 = x[32] & n5654 ;
  assign n32911 = ~n5656 ;
  assign n5657 = n5655 & n32911 ;
  assign n32912 = ~n5450 ;
  assign n5658 = n5447 & n32912 ;
  assign n5659 = n5453 | n5607 ;
  assign n32913 = ~n5658 ;
  assign n5660 = n32913 & n5659 ;
  assign n5661 = n5657 & n5660 ;
  assign n5662 = n5657 | n5660 ;
  assign n32914 = ~n5661 ;
  assign n5663 = n32914 & n5662 ;
  assign n32915 = ~n5601 ;
  assign n5664 = n5462 & n32915 ;
  assign n32916 = ~n5604 ;
  assign n5665 = n5460 & n32916 ;
  assign n5666 = n5664 | n5665 ;
  assign n32917 = ~n5591 ;
  assign n5667 = n32917 & n5598 ;
  assign n5668 = n5590 | n5667 ;
  assign n32918 = ~n5569 ;
  assign n5669 = n5471 & n32918 ;
  assign n5670 = n5568 | n5669 ;
  assign n5671 = n5555 | n5565 ;
  assign n32919 = ~n5504 ;
  assign n5672 = n5488 & n32919 ;
  assign n32920 = ~n5507 ;
  assign n5673 = n32920 & n5514 ;
  assign n5674 = n5672 | n5673 ;
  assign n32921 = ~n5489 ;
  assign n5675 = n5081 & n32921 ;
  assign n32922 = ~n5492 ;
  assign n5676 = n32922 & n5501 ;
  assign n5677 = n5675 | n5676 ;
  assign n27780 = x[87] & n27215 ;
  assign n857 = x[88] & n805 ;
  assign n5678 = n27780 | n857 ;
  assign n32923 = ~n5678 ;
  assign n5679 = x[23] & n32923 ;
  assign n5680 = n28221 & n5678 ;
  assign n5681 = n5679 | n5680 ;
  assign n32924 = ~n5681 ;
  assign n5682 = n5489 & n32924 ;
  assign n5683 = n32921 & n5681 ;
  assign n5684 = n5682 | n5683 ;
  assign n2050 = n1006 & n2046 ;
  assign n911 = x[89] & n900 ;
  assign n965 = x[90] & n949 ;
  assign n5685 = n911 | n965 ;
  assign n5686 = x[91] & n881 ;
  assign n5687 = n5685 | n5686 ;
  assign n5688 = n2050 | n5687 ;
  assign n32925 = ~n5688 ;
  assign n5689 = x[62] & n32925 ;
  assign n5690 = n30886 & n5688 ;
  assign n5691 = n5689 | n5690 ;
  assign n5692 = n5684 | n5691 ;
  assign n5693 = n5684 & n5691 ;
  assign n32926 = ~n5693 ;
  assign n5694 = n5692 & n32926 ;
  assign n32927 = ~n5677 ;
  assign n5695 = n32927 & n5694 ;
  assign n32928 = ~n5694 ;
  assign n5696 = n5677 & n32928 ;
  assign n5697 = n5695 | n5696 ;
  assign n2414 = n1217 & n2410 ;
  assign n1122 = x[92] & n1079 ;
  assign n1166 = x[93] & n1144 ;
  assign n5698 = n1122 | n1166 ;
  assign n5699 = x[94] & n1075 ;
  assign n5700 = n5698 | n5699 ;
  assign n5701 = n2414 | n5700 ;
  assign n32929 = ~n5701 ;
  assign n5702 = x[59] & n32929 ;
  assign n5703 = n30638 & n5701 ;
  assign n5704 = n5702 | n5703 ;
  assign n32930 = ~n5704 ;
  assign n5705 = n5697 & n32930 ;
  assign n32931 = ~n5697 ;
  assign n5706 = n32931 & n5704 ;
  assign n5707 = n5705 | n5706 ;
  assign n32932 = ~n5707 ;
  assign n5708 = n5674 & n32932 ;
  assign n32933 = ~n5674 ;
  assign n5709 = n32933 & n5707 ;
  assign n5710 = n5708 | n5709 ;
  assign n2441 = n1457 & n2438 ;
  assign n1371 = x[95] & n1319 ;
  assign n1419 = x[96] & n1384 ;
  assign n5711 = n1371 | n1419 ;
  assign n5712 = x[97] & n1315 ;
  assign n5713 = n5711 | n5712 ;
  assign n5714 = n2441 | n5713 ;
  assign n32934 = ~n5714 ;
  assign n5715 = x[56] & n32934 ;
  assign n5716 = n30379 & n5714 ;
  assign n5717 = n5715 | n5716 ;
  assign n32935 = ~n5517 ;
  assign n5718 = n32935 & n5518 ;
  assign n32936 = ~n5521 ;
  assign n5719 = n32936 & n5528 ;
  assign n5720 = n5718 | n5719 ;
  assign n5721 = n5717 | n5720 ;
  assign n5722 = n5717 & n5720 ;
  assign n32937 = ~n5722 ;
  assign n5723 = n5721 & n32937 ;
  assign n32938 = ~n5710 ;
  assign n5724 = n32938 & n5723 ;
  assign n32939 = ~n5723 ;
  assign n5725 = n5710 & n32939 ;
  assign n5726 = n5724 | n5725 ;
  assign n2470 = n1690 & n2466 ;
  assign n1602 = x[98] & n1551 ;
  assign n1673 = x[99] & n1616 ;
  assign n5727 = n1602 | n1673 ;
  assign n5728 = x[100] & n1547 ;
  assign n5729 = n5727 | n5728 ;
  assign n5730 = n2470 | n5729 ;
  assign n32940 = ~n5730 ;
  assign n5731 = x[53] & n32940 ;
  assign n5732 = n30125 & n5730 ;
  assign n5733 = n5731 | n5732 ;
  assign n5734 = n5726 | n5733 ;
  assign n5735 = n5726 & n5733 ;
  assign n32941 = ~n5735 ;
  assign n5736 = n5734 & n32941 ;
  assign n32942 = ~n5531 ;
  assign n5737 = n5485 & n32942 ;
  assign n32943 = ~n5534 ;
  assign n5738 = n5482 & n32943 ;
  assign n5739 = n5737 | n5738 ;
  assign n32944 = ~n5739 ;
  assign n5740 = n5736 & n32944 ;
  assign n32945 = ~n5736 ;
  assign n5741 = n32945 & n5739 ;
  assign n5742 = n5740 | n5741 ;
  assign n2631 = n2007 & n2626 ;
  assign n1877 = x[101] & n1866 ;
  assign n1943 = x[102] & n1931 ;
  assign n5743 = n1877 | n1943 ;
  assign n5744 = x[103] & n1862 ;
  assign n5745 = n5743 | n5744 ;
  assign n5746 = n2631 | n5745 ;
  assign n32946 = ~n5746 ;
  assign n5747 = x[50] & n32946 ;
  assign n5748 = n29865 & n5746 ;
  assign n5749 = n5747 | n5748 ;
  assign n5750 = n5742 | n5749 ;
  assign n5751 = n5742 & n5749 ;
  assign n32947 = ~n5751 ;
  assign n5752 = n5750 & n32947 ;
  assign n32948 = ~n5537 ;
  assign n5753 = n5475 & n32948 ;
  assign n32949 = ~n5540 ;
  assign n5754 = n32949 & n5547 ;
  assign n5755 = n5753 | n5754 ;
  assign n32950 = ~n5755 ;
  assign n5756 = n5752 & n32950 ;
  assign n32951 = ~n5752 ;
  assign n5757 = n32951 & n5755 ;
  assign n5758 = n5756 | n5757 ;
  assign n3230 = n2321 & n3223 ;
  assign n2219 = x[104] & n2179 ;
  assign n2290 = x[105] & n2244 ;
  assign n5759 = n2219 | n2290 ;
  assign n5760 = x[106] & n2175 ;
  assign n5761 = n5759 | n5760 ;
  assign n5762 = n3230 | n5761 ;
  assign n32952 = ~n5762 ;
  assign n5763 = x[47] & n32952 ;
  assign n5764 = n29621 & n5762 ;
  assign n5765 = n5763 | n5764 ;
  assign n5766 = n5758 | n5765 ;
  assign n5767 = n5758 & n5765 ;
  assign n32953 = ~n5767 ;
  assign n5768 = n5766 & n32953 ;
  assign n5769 = n5671 & n5768 ;
  assign n5770 = n5671 | n5768 ;
  assign n32954 = ~n5769 ;
  assign n5771 = n32954 & n5770 ;
  assign n3644 = n2635 & n3639 ;
  assign n2526 = x[107] & n2492 ;
  assign n2607 = x[108] & n2557 ;
  assign n5772 = n2526 | n2607 ;
  assign n5773 = x[109] & n2488 ;
  assign n5774 = n5772 | n5773 ;
  assign n5775 = n3644 | n5774 ;
  assign n32955 = ~n5775 ;
  assign n5776 = x[44] & n32955 ;
  assign n5777 = n29400 & n5775 ;
  assign n5778 = n5776 | n5777 ;
  assign n32956 = ~n5778 ;
  assign n5779 = n5771 & n32956 ;
  assign n32957 = ~n5771 ;
  assign n5780 = n32957 & n5778 ;
  assign n5781 = n5779 | n5780 ;
  assign n32958 = ~n5781 ;
  assign n5782 = n5670 & n32958 ;
  assign n32959 = ~n5670 ;
  assign n5783 = n32959 & n5781 ;
  assign n5784 = n5782 | n5783 ;
  assign n4444 = n3162 & n4442 ;
  assign n3060 = x[110] & n3031 ;
  assign n3141 = x[111] & n3096 ;
  assign n5785 = n3060 | n3141 ;
  assign n5786 = x[112] & n3027 ;
  assign n5787 = n5785 | n5786 ;
  assign n5788 = n4444 | n5787 ;
  assign n32960 = ~n5788 ;
  assign n5789 = x[41] & n32960 ;
  assign n5790 = n29184 & n5788 ;
  assign n5791 = n5789 | n5790 ;
  assign n5792 = n5784 | n5791 ;
  assign n5793 = n5784 & n5791 ;
  assign n32961 = ~n5793 ;
  assign n5794 = n5792 & n32961 ;
  assign n32962 = ~n5572 ;
  assign n5795 = n5464 & n32962 ;
  assign n32963 = ~n5575 ;
  assign n5796 = n32963 & n5582 ;
  assign n5797 = n5795 | n5796 ;
  assign n5798 = n5794 | n5797 ;
  assign n5799 = n5794 & n5797 ;
  assign n32964 = ~n5799 ;
  assign n5800 = n5798 & n32964 ;
  assign n4481 = n3574 & n4474 ;
  assign n3456 = x[113] & n3443 ;
  assign n3529 = x[114] & n3508 ;
  assign n5801 = n3456 | n3529 ;
  assign n5802 = x[115] & n3439 ;
  assign n5803 = n5801 | n5802 ;
  assign n5804 = n4481 | n5803 ;
  assign n32965 = ~n5804 ;
  assign n5805 = x[38] & n32965 ;
  assign n5806 = n28996 & n5804 ;
  assign n5807 = n5805 | n5806 ;
  assign n32966 = ~n5800 ;
  assign n5809 = n32966 & n5807 ;
  assign n32967 = ~n5807 ;
  assign n5808 = n5800 & n32967 ;
  assign n32968 = ~n5808 ;
  assign n5810 = n5668 & n32968 ;
  assign n32969 = ~n5809 ;
  assign n5811 = n32969 & n5810 ;
  assign n32970 = ~n5811 ;
  assign n5813 = n5668 & n32970 ;
  assign n5812 = n5809 | n5810 ;
  assign n5814 = n5808 | n5812 ;
  assign n32971 = ~n5813 ;
  assign n5815 = n32971 & n5814 ;
  assign n4059 = n784 & n4041 ;
  assign n3955 = x[116] & n3910 ;
  assign n4014 = x[117] & n3975 ;
  assign n5816 = n3955 | n4014 ;
  assign n5817 = x[118] & n3906 ;
  assign n5818 = n5816 | n5817 ;
  assign n5819 = n4059 | n5818 ;
  assign n32972 = ~n5819 ;
  assign n5820 = x[35] & n32972 ;
  assign n5821 = n28822 & n5819 ;
  assign n5822 = n5820 | n5821 ;
  assign n5823 = n5815 | n5822 ;
  assign n5824 = n5815 & n5822 ;
  assign n32973 = ~n5824 ;
  assign n5825 = n5823 & n32973 ;
  assign n5826 = n5666 | n5825 ;
  assign n5827 = n5666 & n5825 ;
  assign n32974 = ~n5827 ;
  assign n5828 = n5826 & n32974 ;
  assign n5829 = n5663 | n5828 ;
  assign n5860 = n5663 & n5828 ;
  assign n32975 = ~n5860 ;
  assign n5861 = n5859 & n32975 ;
  assign n5862 = n5829 & n5861 ;
  assign n32976 = ~n5862 ;
  assign n5863 = n5859 & n32976 ;
  assign n5864 = n5860 | n5862 ;
  assign n32977 = ~n5864 ;
  assign n5865 = n5829 & n32977 ;
  assign n5866 = n5863 | n5865 ;
  assign n32978 = ~n5866 ;
  assign n5868 = n5650 & n32978 ;
  assign n32979 = ~n5650 ;
  assign n5869 = n32979 & n5866 ;
  assign n5870 = n5868 | n5869 ;
  assign n32980 = ~n5870 ;
  assign n23195 = n5619 & n32980 ;
  assign n32981 = ~n5619 ;
  assign n23196 = n32981 & n5870 ;
  assign n23197 = n23195 | n23196 ;
  assign n23198 = n23194 & n23197 ;
  assign n27781 = n23194 | n23196 ;
  assign n27782 = n23195 | n27781 ;
  assign n32982 = ~n23198 ;
  assign n216 = n32982 & n27782 ;
  assign n5871 = n5619 & n5870 ;
  assign n23199 = n5871 | n23198 ;
  assign n5867 = n5650 & n5866 ;
  assign n23200 = n5649 | n5867 ;
  assign n4641 = n642 & n4632 ;
  assign n4533 = x[123] & n4514 ;
  assign n4622 = x[124] & n4572 ;
  assign n23201 = n4533 | n4622 ;
  assign n23202 = x[125] & n4504 ;
  assign n23203 = n23201 | n23202 ;
  assign n23204 = n4641 | n23203 ;
  assign n32983 = ~n23204 ;
  assign n23205 = x[29] & n32983 ;
  assign n23206 = n28483 & n23204 ;
  assign n23207 = n23205 | n23206 ;
  assign n32984 = ~n5660 ;
  assign n23208 = n5657 & n32984 ;
  assign n32985 = ~n23208 ;
  assign n23209 = n5829 & n32985 ;
  assign n23210 = n23207 & n23209 ;
  assign n23211 = n23207 | n23209 ;
  assign n32986 = ~n23210 ;
  assign n23212 = n32986 & n23211 ;
  assign n32987 = ~n5815 ;
  assign n23213 = n32987 & n5822 ;
  assign n32988 = ~n5825 ;
  assign n23214 = n5666 & n32988 ;
  assign n23215 = n23213 | n23214 ;
  assign n659 = x[122] & n652 ;
  assign n23216 = x[120] & n663 ;
  assign n23217 = x[121] & n720 ;
  assign n23218 = n23216 | n23217 ;
  assign n23219 = n659 | n23218 ;
  assign n23220 = n779 & n5022 ;
  assign n23221 = n23219 | n23220 ;
  assign n23222 = n28658 & n23221 ;
  assign n32989 = ~n23221 ;
  assign n23223 = x[32] & n32989 ;
  assign n23224 = n23222 | n23223 ;
  assign n32990 = ~n23224 ;
  assign n23225 = n23215 & n32990 ;
  assign n32991 = ~n23215 ;
  assign n23226 = n32991 & n23224 ;
  assign n23227 = n23225 | n23226 ;
  assign n32992 = ~n5742 ;
  assign n23228 = n32992 & n5749 ;
  assign n23229 = n5757 | n23228 ;
  assign n3007 = n2007 & n3001 ;
  assign n1887 = x[102] & n1866 ;
  assign n1948 = x[103] & n1931 ;
  assign n23294 = n1887 | n1948 ;
  assign n23295 = x[104] & n1862 ;
  assign n23296 = n23294 | n23295 ;
  assign n23297 = n3007 | n23296 ;
  assign n23298 = x[50] | n23297 ;
  assign n23299 = x[50] & n23297 ;
  assign n32993 = ~n23299 ;
  assign n23300 = n23298 & n32993 ;
  assign n32994 = ~n5726 ;
  assign n23230 = n32994 & n5733 ;
  assign n23231 = n5741 | n23230 ;
  assign n32995 = ~n5684 ;
  assign n23232 = n32995 & n5691 ;
  assign n23233 = n5696 | n23232 ;
  assign n279 = x[88] & n27215 ;
  assign n858 = x[89] & n805 ;
  assign n23234 = n279 | n858 ;
  assign n23235 = n5680 | n5682 ;
  assign n32996 = ~n23235 ;
  assign n23236 = n23234 & n32996 ;
  assign n32997 = ~n23234 ;
  assign n23237 = n32997 & n23235 ;
  assign n23238 = n23236 | n23237 ;
  assign n886 = x[92] & n881 ;
  assign n23239 = x[90] & n900 ;
  assign n23240 = x[91] & n949 ;
  assign n23241 = n23239 | n23240 ;
  assign n23242 = n886 | n23241 ;
  assign n23243 = n1006 & n1841 ;
  assign n23244 = n23242 | n23243 ;
  assign n23245 = n30886 & n23244 ;
  assign n32998 = ~n23244 ;
  assign n23246 = x[62] & n32998 ;
  assign n23247 = n23245 | n23246 ;
  assign n32999 = ~n23247 ;
  assign n23248 = n23238 & n32999 ;
  assign n33000 = ~n23238 ;
  assign n23249 = n33000 & n23247 ;
  assign n23250 = n23248 | n23249 ;
  assign n33001 = ~n23250 ;
  assign n23251 = n23233 & n33001 ;
  assign n33002 = ~n23233 ;
  assign n23252 = n33002 & n23250 ;
  assign n23253 = n23251 | n23252 ;
  assign n2159 = n1217 & n2152 ;
  assign n1104 = x[93] & n1079 ;
  assign n1180 = x[94] & n1144 ;
  assign n23254 = n1104 | n1180 ;
  assign n23255 = x[95] & n1075 ;
  assign n23256 = n23254 | n23255 ;
  assign n23257 = n2159 | n23256 ;
  assign n33003 = ~n23257 ;
  assign n23258 = x[59] & n33003 ;
  assign n23259 = n30638 & n23257 ;
  assign n23260 = n23258 | n23259 ;
  assign n23261 = n23253 | n23260 ;
  assign n23262 = n23253 & n23260 ;
  assign n33004 = ~n23262 ;
  assign n23263 = n23261 & n33004 ;
  assign n23264 = n5706 | n5708 ;
  assign n33005 = ~n23264 ;
  assign n23265 = n23263 & n33005 ;
  assign n33006 = ~n23263 ;
  assign n23266 = n33006 & n23264 ;
  assign n23267 = n23265 | n23266 ;
  assign n2848 = n1457 & n2841 ;
  assign n1359 = x[96] & n1319 ;
  assign n1405 = x[97] & n1384 ;
  assign n23268 = n1359 | n1405 ;
  assign n23269 = x[98] & n1315 ;
  assign n23270 = n23268 | n23269 ;
  assign n23271 = n2848 | n23270 ;
  assign n33007 = ~n23271 ;
  assign n23272 = x[56] & n33007 ;
  assign n23273 = n30379 & n23271 ;
  assign n23274 = n23272 | n23273 ;
  assign n23275 = n23267 | n23274 ;
  assign n23276 = n23267 & n23274 ;
  assign n33008 = ~n23276 ;
  assign n23277 = n23275 & n33008 ;
  assign n23278 = n5722 | n5724 ;
  assign n23279 = n23277 | n23278 ;
  assign n23280 = n23277 & n23278 ;
  assign n33009 = ~n23280 ;
  assign n23281 = n23279 & n33009 ;
  assign n2983 = n1690 & n2977 ;
  assign n1571 = x[99] & n1551 ;
  assign n1656 = x[100] & n1616 ;
  assign n23282 = n1571 | n1656 ;
  assign n23283 = x[101] & n1547 ;
  assign n23284 = n23282 | n23283 ;
  assign n23285 = n2983 | n23284 ;
  assign n33010 = ~n23285 ;
  assign n23286 = x[53] & n33010 ;
  assign n23287 = n30125 & n23285 ;
  assign n23288 = n23286 | n23287 ;
  assign n23289 = n23281 | n23288 ;
  assign n23290 = n23281 & n23288 ;
  assign n33011 = ~n23290 ;
  assign n23291 = n23289 & n33011 ;
  assign n23292 = n23231 | n23291 ;
  assign n23293 = n23231 & n23291 ;
  assign n33012 = ~n23293 ;
  assign n23301 = n23292 & n33012 ;
  assign n33013 = ~n23301 ;
  assign n23302 = n23300 & n33013 ;
  assign n33014 = ~n23300 ;
  assign n23303 = n23292 & n33014 ;
  assign n23304 = n33012 & n23303 ;
  assign n23305 = n23302 | n23304 ;
  assign n33015 = ~n23229 ;
  assign n23306 = n33015 & n23305 ;
  assign n33016 = ~n23305 ;
  assign n23307 = n23229 & n33016 ;
  assign n23308 = n23306 | n23307 ;
  assign n3206 = n2321 & n3199 ;
  assign n2185 = x[105] & n2179 ;
  assign n2275 = x[106] & n2244 ;
  assign n23309 = n2185 | n2275 ;
  assign n23310 = x[107] & n2175 ;
  assign n23311 = n23309 | n23310 ;
  assign n23312 = n3206 | n23311 ;
  assign n33017 = ~n23312 ;
  assign n23313 = x[47] & n33017 ;
  assign n23314 = n29621 & n23312 ;
  assign n23315 = n23313 | n23314 ;
  assign n23316 = n23308 | n23315 ;
  assign n23317 = n23308 & n23315 ;
  assign n33018 = ~n23317 ;
  assign n23318 = n23316 & n33018 ;
  assign n33019 = ~n5758 ;
  assign n23319 = n33019 & n5765 ;
  assign n33020 = ~n5768 ;
  assign n23320 = n5671 & n33020 ;
  assign n23321 = n23319 | n23320 ;
  assign n23322 = n23318 | n23321 ;
  assign n23323 = n23318 & n23321 ;
  assign n33021 = ~n23323 ;
  assign n23324 = n23322 & n33021 ;
  assign n3616 = n2635 & n3615 ;
  assign n2539 = x[108] & n2492 ;
  assign n2575 = x[109] & n2557 ;
  assign n23325 = n2539 | n2575 ;
  assign n23326 = x[110] & n2488 ;
  assign n23327 = n23325 | n23326 ;
  assign n23328 = n3616 | n23327 ;
  assign n33022 = ~n23328 ;
  assign n23329 = x[44] & n33022 ;
  assign n23330 = n29400 & n23328 ;
  assign n23331 = n23329 | n23330 ;
  assign n23332 = n23324 | n23331 ;
  assign n23333 = n23324 & n23331 ;
  assign n33023 = ~n23333 ;
  assign n23334 = n23332 & n33023 ;
  assign n23335 = n5780 | n5782 ;
  assign n33024 = ~n23335 ;
  assign n23336 = n23334 & n33024 ;
  assign n33025 = ~n23334 ;
  assign n23337 = n33025 & n23335 ;
  assign n23338 = n23336 | n23337 ;
  assign n4094 = n3162 & n4087 ;
  assign n3041 = x[111] & n3031 ;
  assign n3112 = x[112] & n3096 ;
  assign n23339 = n3041 | n3112 ;
  assign n23340 = x[113] & n3027 ;
  assign n23341 = n23339 | n23340 ;
  assign n23342 = n4094 | n23341 ;
  assign n33026 = ~n23342 ;
  assign n23343 = x[41] & n33026 ;
  assign n23344 = n29184 & n23342 ;
  assign n23345 = n23343 | n23344 ;
  assign n23346 = n23338 | n23345 ;
  assign n23347 = n23338 & n23345 ;
  assign n33027 = ~n23347 ;
  assign n23348 = n23346 & n33027 ;
  assign n33028 = ~n5784 ;
  assign n23349 = n33028 & n5791 ;
  assign n33029 = ~n5794 ;
  assign n23350 = n33029 & n5797 ;
  assign n23351 = n23349 | n23350 ;
  assign n33030 = ~n23351 ;
  assign n23352 = n23348 & n33030 ;
  assign n33031 = ~n23348 ;
  assign n23353 = n33031 & n23351 ;
  assign n23354 = n23352 | n23353 ;
  assign n4703 = n3574 & n4702 ;
  assign n3449 = x[114] & n3443 ;
  assign n3565 = x[115] & n3508 ;
  assign n23355 = n3449 | n3565 ;
  assign n23356 = x[116] & n3439 ;
  assign n23357 = n23355 | n23356 ;
  assign n23358 = n4703 | n23357 ;
  assign n33032 = ~n23358 ;
  assign n23359 = x[38] & n33032 ;
  assign n23360 = n28996 & n23358 ;
  assign n23361 = n23359 | n23360 ;
  assign n23362 = n23354 | n23361 ;
  assign n23363 = n23354 & n23361 ;
  assign n33033 = ~n23363 ;
  assign n23364 = n23362 & n33033 ;
  assign n23365 = n5812 & n23364 ;
  assign n23366 = n5812 | n23364 ;
  assign n33034 = ~n23365 ;
  assign n23367 = n33034 & n23366 ;
  assign n5048 = n4041 & n5047 ;
  assign n3914 = x[117] & n3910 ;
  assign n4008 = x[118] & n3975 ;
  assign n23368 = n3914 | n4008 ;
  assign n23369 = x[119] & n3906 ;
  assign n23370 = n23368 | n23369 ;
  assign n23371 = n5048 | n23370 ;
  assign n33035 = ~n23371 ;
  assign n23372 = x[35] & n33035 ;
  assign n23373 = n28822 & n23371 ;
  assign n23374 = n23372 | n23373 ;
  assign n33036 = ~n23374 ;
  assign n23375 = n23367 & n33036 ;
  assign n33037 = ~n23367 ;
  assign n23376 = n33037 & n23374 ;
  assign n23377 = n23375 | n23376 ;
  assign n33038 = ~n23377 ;
  assign n23378 = n23227 & n33038 ;
  assign n33039 = ~n23227 ;
  assign n23379 = n33039 & n23377 ;
  assign n23380 = n23378 | n23379 ;
  assign n33040 = ~n23380 ;
  assign n23381 = n23212 & n33040 ;
  assign n33041 = ~n23212 ;
  assign n23382 = n33041 & n23380 ;
  assign n23383 = n23381 | n23382 ;
  assign n23384 = n5858 | n5862 ;
  assign n6191 = n452 & n6186 ;
  assign n23385 = x[126] & n330 ;
  assign n23386 = x[127] & n390 ;
  assign n23387 = n23385 | n23386 ;
  assign n23388 = n6191 | n23387 ;
  assign n33042 = ~n23388 ;
  assign n23389 = x[26] & n33042 ;
  assign n23390 = n28342 & n23388 ;
  assign n23391 = n23389 | n23390 ;
  assign n33043 = ~n23391 ;
  assign n23392 = n23384 & n33043 ;
  assign n33044 = ~n23384 ;
  assign n23393 = n33044 & n23391 ;
  assign n23394 = n23392 | n23393 ;
  assign n23396 = n23383 & n23394 ;
  assign n23395 = n23383 | n23393 ;
  assign n23397 = n23392 | n23395 ;
  assign n33045 = ~n23396 ;
  assign n23398 = n33045 & n23397 ;
  assign n33046 = ~n23398 ;
  assign n23399 = n23200 & n33046 ;
  assign n33047 = ~n23200 ;
  assign n23400 = n33047 & n23398 ;
  assign n23401 = n23399 | n23400 ;
  assign n23402 = n23199 & n23401 ;
  assign n23403 = n23199 | n23400 ;
  assign n23404 = n23399 | n23403 ;
  assign n33048 = ~n23402 ;
  assign n217 = n33048 & n23404 ;
  assign n23406 = n23200 & n23398 ;
  assign n23407 = n23402 | n23406 ;
  assign n23408 = n23384 & n23391 ;
  assign n23409 = n23396 | n23408 ;
  assign n33049 = ~n23209 ;
  assign n23410 = n23207 & n33049 ;
  assign n23411 = n23212 | n23380 ;
  assign n33050 = ~n23410 ;
  assign n23412 = n33050 & n23411 ;
  assign n389 = x[127] & n330 ;
  assign n5361 = n452 & n5360 ;
  assign n23413 = n389 | n5361 ;
  assign n33051 = ~n23413 ;
  assign n23414 = x[26] & n33051 ;
  assign n23415 = n28342 & n23413 ;
  assign n23416 = n23414 | n23415 ;
  assign n33052 = ~n23416 ;
  assign n23417 = n23412 & n33052 ;
  assign n33053 = ~n23412 ;
  assign n23418 = n33053 & n23416 ;
  assign n23419 = n23417 | n23418 ;
  assign n5397 = n4632 & n5388 ;
  assign n4570 = x[124] & n4514 ;
  assign n4626 = x[125] & n4572 ;
  assign n23420 = n4570 | n4626 ;
  assign n23421 = x[126] & n4504 ;
  assign n23422 = n23420 | n23421 ;
  assign n23423 = n5397 | n23422 ;
  assign n33054 = ~n23423 ;
  assign n23424 = x[29] & n33054 ;
  assign n23425 = n28483 & n23423 ;
  assign n23426 = n23424 | n23425 ;
  assign n23427 = n23215 & n23224 ;
  assign n23428 = n23378 | n23427 ;
  assign n23429 = n23426 | n23428 ;
  assign n23430 = n23426 & n23428 ;
  assign n33055 = ~n23430 ;
  assign n23431 = n23429 & n33055 ;
  assign n5426 = n779 & n5417 ;
  assign n673 = x[121] & n663 ;
  assign n774 = x[122] & n720 ;
  assign n23432 = n673 | n774 ;
  assign n23433 = x[123] & n652 ;
  assign n23434 = n23432 | n23433 ;
  assign n23435 = n5426 | n23434 ;
  assign n23436 = x[32] | n23435 ;
  assign n23437 = x[32] & n23435 ;
  assign n33056 = ~n23437 ;
  assign n23438 = n23436 & n33056 ;
  assign n33057 = ~n23364 ;
  assign n23439 = n5812 & n33057 ;
  assign n23440 = n23376 | n23439 ;
  assign n33058 = ~n23440 ;
  assign n23441 = n23438 & n33058 ;
  assign n33059 = ~n23438 ;
  assign n23442 = n33059 & n23440 ;
  assign n23443 = n23441 | n23442 ;
  assign n4682 = n4041 & n4678 ;
  assign n3922 = x[118] & n3910 ;
  assign n3995 = x[119] & n3975 ;
  assign n23444 = n3922 | n3995 ;
  assign n23445 = x[120] & n3906 ;
  assign n23446 = n23444 | n23445 ;
  assign n23447 = n4682 | n23446 ;
  assign n33060 = ~n23447 ;
  assign n23448 = x[35] & n33060 ;
  assign n23449 = n28822 & n23447 ;
  assign n23450 = n23448 | n23449 ;
  assign n33061 = ~n23354 ;
  assign n23451 = n33061 & n23361 ;
  assign n23452 = n23353 | n23451 ;
  assign n3577 = n797 & n3574 ;
  assign n3447 = x[115] & n3443 ;
  assign n3563 = x[116] & n3508 ;
  assign n23579 = n3447 | n3563 ;
  assign n23580 = x[117] & n3439 ;
  assign n23581 = n23579 | n23580 ;
  assign n23582 = n3577 | n23581 ;
  assign n23583 = x[38] | n23582 ;
  assign n23584 = x[38] & n23582 ;
  assign n33062 = ~n23584 ;
  assign n23585 = n23583 & n33062 ;
  assign n33063 = ~n23338 ;
  assign n23453 = n33063 & n23345 ;
  assign n23454 = n23337 | n23453 ;
  assign n33064 = ~n23308 ;
  assign n23455 = n33064 & n23315 ;
  assign n23456 = n23307 | n23455 ;
  assign n3881 = n2321 & n3876 ;
  assign n2214 = x[106] & n2179 ;
  assign n2259 = x[107] & n2244 ;
  assign n23457 = n2214 | n2259 ;
  assign n23458 = x[108] & n2175 ;
  assign n23459 = n23457 | n23458 ;
  assign n23460 = n3881 | n23459 ;
  assign n33065 = ~n23460 ;
  assign n23461 = x[47] & n33065 ;
  assign n23462 = n29621 & n23460 ;
  assign n23463 = n23461 | n23462 ;
  assign n33066 = ~n23291 ;
  assign n23464 = n23231 & n33066 ;
  assign n23465 = n23302 | n23464 ;
  assign n33067 = ~n23267 ;
  assign n23466 = n33067 & n23274 ;
  assign n23467 = n23266 | n23466 ;
  assign n2317 = n1457 & n2313 ;
  assign n1343 = x[97] & n1319 ;
  assign n1412 = x[98] & n1384 ;
  assign n23468 = n1343 | n1412 ;
  assign n23469 = x[99] & n1315 ;
  assign n23470 = n23468 | n23469 ;
  assign n23471 = n2317 | n23470 ;
  assign n33068 = ~n23471 ;
  assign n23472 = x[56] & n33068 ;
  assign n23473 = n30379 & n23471 ;
  assign n23474 = n23472 | n23473 ;
  assign n33069 = ~n23253 ;
  assign n23475 = n33069 & n23260 ;
  assign n23476 = n23251 | n23475 ;
  assign n2004 = n1217 & n2000 ;
  assign n1127 = x[94] & n1079 ;
  assign n1184 = x[95] & n1144 ;
  assign n23477 = n1127 | n1184 ;
  assign n23478 = x[96] & n1075 ;
  assign n23479 = n23477 | n23478 ;
  assign n23480 = n2004 | n23479 ;
  assign n23481 = x[59] | n23480 ;
  assign n23482 = x[59] & n23480 ;
  assign n33070 = ~n23482 ;
  assign n23483 = n23481 & n33070 ;
  assign n23484 = n23237 | n23249 ;
  assign n280 = x[89] & n27215 ;
  assign n861 = x[90] & n805 ;
  assign n23485 = n280 | n861 ;
  assign n23486 = n23234 | n23485 ;
  assign n23487 = n23234 & n23485 ;
  assign n33071 = ~n23487 ;
  assign n23488 = n23486 & n33071 ;
  assign n884 = x[93] & n881 ;
  assign n23489 = x[91] & n900 ;
  assign n23490 = x[92] & n949 ;
  assign n23491 = n23489 | n23490 ;
  assign n23492 = n884 | n23491 ;
  assign n23493 = n1006 & n1685 ;
  assign n23494 = n23492 | n23493 ;
  assign n23495 = n30886 & n23494 ;
  assign n33072 = ~n23494 ;
  assign n23496 = x[62] & n33072 ;
  assign n23497 = n23495 | n23496 ;
  assign n23498 = n23488 | n23497 ;
  assign n23499 = n23488 & n23497 ;
  assign n33073 = ~n23499 ;
  assign n23500 = n23498 & n33073 ;
  assign n33074 = ~n23500 ;
  assign n23501 = n23484 & n33074 ;
  assign n33075 = ~n23484 ;
  assign n23502 = n33075 & n23500 ;
  assign n23503 = n23501 | n23502 ;
  assign n33076 = ~n23503 ;
  assign n23504 = n23483 & n33076 ;
  assign n33077 = ~n23483 ;
  assign n23505 = n33077 & n23503 ;
  assign n23506 = n23504 | n23505 ;
  assign n23507 = n23476 | n23506 ;
  assign n23508 = n23476 & n23506 ;
  assign n33078 = ~n23508 ;
  assign n23509 = n23507 & n33078 ;
  assign n23510 = n23474 | n23509 ;
  assign n23511 = n23474 & n23509 ;
  assign n33079 = ~n23511 ;
  assign n23512 = n23510 & n33079 ;
  assign n23513 = n23467 | n23512 ;
  assign n23514 = n23467 & n23512 ;
  assign n33080 = ~n23514 ;
  assign n23515 = n23513 & n33080 ;
  assign n2873 = n1690 & n2867 ;
  assign n1573 = x[100] & n1551 ;
  assign n1639 = x[101] & n1616 ;
  assign n23516 = n1573 | n1639 ;
  assign n23517 = x[102] & n1547 ;
  assign n23518 = n23516 | n23517 ;
  assign n23519 = n2873 | n23518 ;
  assign n33081 = ~n23519 ;
  assign n23520 = x[53] & n33081 ;
  assign n23521 = n30125 & n23519 ;
  assign n23522 = n23520 | n23521 ;
  assign n23523 = n23515 | n23522 ;
  assign n23524 = n23515 & n23522 ;
  assign n33082 = ~n23524 ;
  assign n23525 = n23523 & n33082 ;
  assign n33083 = ~n23277 ;
  assign n23526 = n33083 & n23278 ;
  assign n33084 = ~n23281 ;
  assign n23527 = n33084 & n23288 ;
  assign n23528 = n23526 | n23527 ;
  assign n33085 = ~n23528 ;
  assign n23529 = n23525 & n33085 ;
  assign n33086 = ~n23525 ;
  assign n23530 = n33086 & n23528 ;
  assign n23531 = n23529 | n23530 ;
  assign n3415 = n2007 & n3409 ;
  assign n1886 = x[103] & n1866 ;
  assign n1958 = x[104] & n1931 ;
  assign n23532 = n1886 | n1958 ;
  assign n23533 = x[105] & n1862 ;
  assign n23534 = n23532 | n23533 ;
  assign n23535 = n3415 | n23534 ;
  assign n33087 = ~n23535 ;
  assign n23536 = x[50] & n33087 ;
  assign n23537 = n29865 & n23535 ;
  assign n23538 = n23536 | n23537 ;
  assign n33088 = ~n23538 ;
  assign n23539 = n23531 & n33088 ;
  assign n33089 = ~n23531 ;
  assign n23540 = n33089 & n23538 ;
  assign n23541 = n23539 | n23540 ;
  assign n33090 = ~n23465 ;
  assign n23542 = n33090 & n23541 ;
  assign n33091 = ~n23541 ;
  assign n23543 = n23465 & n33091 ;
  assign n23544 = n23542 | n23543 ;
  assign n23545 = n23463 | n23544 ;
  assign n23546 = n23463 & n23544 ;
  assign n33092 = ~n23546 ;
  assign n23547 = n23545 & n33092 ;
  assign n23548 = n23456 | n23547 ;
  assign n23549 = n23456 & n23547 ;
  assign n33093 = ~n23549 ;
  assign n23550 = n23548 & n33093 ;
  assign n4253 = n2635 & n4246 ;
  assign n2533 = x[109] & n2492 ;
  assign n2568 = x[110] & n2557 ;
  assign n23551 = n2533 | n2568 ;
  assign n23552 = x[111] & n2488 ;
  assign n23553 = n23551 | n23552 ;
  assign n23554 = n4253 | n23553 ;
  assign n33094 = ~n23554 ;
  assign n23555 = x[44] & n33094 ;
  assign n23556 = n29400 & n23554 ;
  assign n23557 = n23555 | n23556 ;
  assign n23558 = n23550 | n23557 ;
  assign n23559 = n23550 & n23557 ;
  assign n33095 = ~n23559 ;
  assign n23560 = n23558 & n33095 ;
  assign n33096 = ~n23318 ;
  assign n23561 = n33096 & n23321 ;
  assign n33097 = ~n23324 ;
  assign n23562 = n33097 & n23331 ;
  assign n23563 = n23561 | n23562 ;
  assign n33098 = ~n23563 ;
  assign n23564 = n23560 & n33098 ;
  assign n33099 = ~n23560 ;
  assign n23565 = n33099 & n23563 ;
  assign n23566 = n23564 | n23565 ;
  assign n4277 = n3162 & n4276 ;
  assign n3055 = x[112] & n3031 ;
  assign n3109 = x[113] & n3096 ;
  assign n23567 = n3055 | n3109 ;
  assign n23568 = x[114] & n3027 ;
  assign n23569 = n23567 | n23568 ;
  assign n23570 = n4277 | n23569 ;
  assign n33100 = ~n23570 ;
  assign n23571 = x[41] & n33100 ;
  assign n23572 = n29184 & n23570 ;
  assign n23573 = n23571 | n23572 ;
  assign n23574 = n23566 | n23573 ;
  assign n23575 = n23566 & n23573 ;
  assign n33101 = ~n23575 ;
  assign n23576 = n23574 & n33101 ;
  assign n23577 = n23454 | n23576 ;
  assign n23578 = n23454 & n23576 ;
  assign n33102 = ~n23578 ;
  assign n23586 = n23577 & n33102 ;
  assign n33103 = ~n23586 ;
  assign n23587 = n23585 & n33103 ;
  assign n33104 = ~n23585 ;
  assign n23588 = n23577 & n33104 ;
  assign n23589 = n33102 & n23588 ;
  assign n23590 = n23587 | n23589 ;
  assign n33105 = ~n23452 ;
  assign n23591 = n33105 & n23590 ;
  assign n33106 = ~n23590 ;
  assign n23592 = n23452 & n33106 ;
  assign n23593 = n23591 | n23592 ;
  assign n23594 = n23450 | n23593 ;
  assign n23595 = n23450 & n23593 ;
  assign n33107 = ~n23595 ;
  assign n23596 = n23594 & n33107 ;
  assign n23597 = n23443 & n23596 ;
  assign n23598 = n23443 | n23596 ;
  assign n33108 = ~n23597 ;
  assign n23599 = n33108 & n23598 ;
  assign n23600 = n23431 & n23599 ;
  assign n23601 = n23431 | n23599 ;
  assign n33109 = ~n23600 ;
  assign n23602 = n33109 & n23601 ;
  assign n33110 = ~n23602 ;
  assign n23603 = n23419 & n33110 ;
  assign n33111 = ~n23419 ;
  assign n23604 = n33111 & n23602 ;
  assign n23605 = n23603 | n23604 ;
  assign n33112 = ~n23409 ;
  assign n23606 = n33112 & n23605 ;
  assign n33113 = ~n23605 ;
  assign n23607 = n23409 & n33113 ;
  assign n23608 = n23606 | n23607 ;
  assign n23609 = n23407 | n23608 ;
  assign n23610 = n23407 & n23608 ;
  assign n33114 = ~n23610 ;
  assign n218 = n23609 & n33114 ;
  assign n23612 = n23419 | n23602 ;
  assign n33115 = ~n23418 ;
  assign n23613 = n33115 & n23612 ;
  assign n33116 = ~n23599 ;
  assign n23614 = n23431 & n33116 ;
  assign n23615 = n23430 | n23614 ;
  assign n5633 = n4632 & n5629 ;
  assign n4568 = x[125] & n4514 ;
  assign n4605 = x[126] & n4572 ;
  assign n23616 = n4568 | n4605 ;
  assign n23617 = x[127] & n4504 ;
  assign n23618 = n23616 | n23617 ;
  assign n23619 = n5633 | n23618 ;
  assign n33117 = ~n23619 ;
  assign n23620 = x[29] & n33117 ;
  assign n23621 = n28483 & n23619 ;
  assign n23622 = n23620 | n23621 ;
  assign n33118 = ~n23622 ;
  assign n23623 = n23615 & n33118 ;
  assign n33119 = ~n23615 ;
  assign n23624 = n33119 & n23622 ;
  assign n23625 = n23623 | n23624 ;
  assign n33120 = ~n23576 ;
  assign n23626 = n23454 & n33120 ;
  assign n23627 = n23587 | n23626 ;
  assign n33121 = ~n23566 ;
  assign n23628 = n33121 & n23573 ;
  assign n23629 = n23565 | n23628 ;
  assign n33122 = ~n23544 ;
  assign n23630 = n23463 & n33122 ;
  assign n23631 = n23543 | n23630 ;
  assign n23632 = n23530 | n23540 ;
  assign n2446 = n1217 & n2438 ;
  assign n1103 = x[95] & n1079 ;
  assign n1167 = x[96] & n1144 ;
  assign n23633 = n1103 | n1167 ;
  assign n23634 = x[97] & n1075 ;
  assign n23635 = n23633 | n23634 ;
  assign n23636 = n2446 | n23635 ;
  assign n23637 = x[59] | n23636 ;
  assign n23638 = x[59] & n23636 ;
  assign n33123 = ~n23638 ;
  assign n23639 = n23637 & n33123 ;
  assign n23640 = n23501 | n23504 ;
  assign n33124 = ~n23640 ;
  assign n23641 = n23639 & n33124 ;
  assign n33125 = ~n23639 ;
  assign n23642 = n33125 & n23640 ;
  assign n23643 = n23641 | n23642 ;
  assign n33126 = ~n23485 ;
  assign n23644 = n23234 & n33126 ;
  assign n33127 = ~n23488 ;
  assign n23645 = n33127 & n23497 ;
  assign n23646 = n23644 | n23645 ;
  assign n281 = x[90] & n27215 ;
  assign n846 = x[91] & n805 ;
  assign n23647 = n281 | n846 ;
  assign n33128 = ~n23647 ;
  assign n23648 = x[26] & n33128 ;
  assign n23649 = n28342 & n23647 ;
  assign n23650 = n23648 | n23649 ;
  assign n33129 = ~n23650 ;
  assign n23651 = n23485 & n33129 ;
  assign n23652 = n33126 & n23650 ;
  assign n23653 = n23651 | n23652 ;
  assign n33130 = ~n23653 ;
  assign n23654 = n23646 & n33130 ;
  assign n33131 = ~n23646 ;
  assign n23655 = n33131 & n23653 ;
  assign n23656 = n23654 | n23655 ;
  assign n2418 = n1006 & n2410 ;
  assign n918 = x[92] & n900 ;
  assign n961 = x[93] & n949 ;
  assign n23657 = n918 | n961 ;
  assign n23658 = x[94] & n881 ;
  assign n23659 = n23657 | n23658 ;
  assign n23660 = n2418 | n23659 ;
  assign n33132 = ~n23660 ;
  assign n23661 = x[62] & n33132 ;
  assign n23662 = n30886 & n23660 ;
  assign n23663 = n23661 | n23662 ;
  assign n23664 = n23656 | n23663 ;
  assign n23665 = n23656 & n23663 ;
  assign n33133 = ~n23665 ;
  assign n23666 = n23664 & n33133 ;
  assign n23667 = n23643 & n23666 ;
  assign n23668 = n23643 | n23666 ;
  assign n33134 = ~n23667 ;
  assign n23669 = n33134 & n23668 ;
  assign n2469 = n1457 & n2466 ;
  assign n1337 = x[98] & n1319 ;
  assign n1398 = x[99] & n1384 ;
  assign n23670 = n1337 | n1398 ;
  assign n23671 = x[100] & n1315 ;
  assign n23672 = n23670 | n23671 ;
  assign n23673 = n2469 | n23672 ;
  assign n33135 = ~n23673 ;
  assign n23674 = x[56] & n33135 ;
  assign n23675 = n30379 & n23673 ;
  assign n23676 = n23674 | n23675 ;
  assign n23677 = n23669 | n23676 ;
  assign n23678 = n23669 & n23676 ;
  assign n33136 = ~n23678 ;
  assign n23679 = n23677 & n33136 ;
  assign n33137 = ~n23506 ;
  assign n23680 = n23476 & n33137 ;
  assign n33138 = ~n23509 ;
  assign n23681 = n23474 & n33138 ;
  assign n23682 = n23680 | n23681 ;
  assign n33139 = ~n23682 ;
  assign n23683 = n23679 & n33139 ;
  assign n33140 = ~n23679 ;
  assign n23684 = n33140 & n23682 ;
  assign n23685 = n23683 | n23684 ;
  assign n2633 = n1690 & n2626 ;
  assign n1570 = x[101] & n1551 ;
  assign n1633 = x[102] & n1616 ;
  assign n23686 = n1570 | n1633 ;
  assign n23687 = x[103] & n1547 ;
  assign n23688 = n23686 | n23687 ;
  assign n23689 = n2633 | n23688 ;
  assign n33141 = ~n23689 ;
  assign n23690 = x[53] & n33141 ;
  assign n23691 = n30125 & n23689 ;
  assign n23692 = n23690 | n23691 ;
  assign n23693 = n23685 | n23692 ;
  assign n23694 = n23685 & n23692 ;
  assign n33142 = ~n23694 ;
  assign n23695 = n23693 & n33142 ;
  assign n33143 = ~n23512 ;
  assign n23696 = n23467 & n33143 ;
  assign n33144 = ~n23515 ;
  assign n23697 = n33144 & n23522 ;
  assign n23698 = n23696 | n23697 ;
  assign n33145 = ~n23698 ;
  assign n23699 = n23695 & n33145 ;
  assign n33146 = ~n23695 ;
  assign n23700 = n33146 & n23698 ;
  assign n23701 = n23699 | n23700 ;
  assign n3232 = n2007 & n3223 ;
  assign n1888 = x[104] & n1866 ;
  assign n1960 = x[105] & n1931 ;
  assign n23702 = n1888 | n1960 ;
  assign n23703 = x[106] & n1862 ;
  assign n23704 = n23702 | n23703 ;
  assign n23705 = n3232 | n23704 ;
  assign n33147 = ~n23705 ;
  assign n23706 = x[50] & n33147 ;
  assign n23707 = n29865 & n23705 ;
  assign n23708 = n23706 | n23707 ;
  assign n23709 = n23701 | n23708 ;
  assign n23710 = n23701 & n23708 ;
  assign n33148 = ~n23710 ;
  assign n23711 = n23709 & n33148 ;
  assign n23712 = n23632 & n23711 ;
  assign n23713 = n23632 | n23711 ;
  assign n33149 = ~n23712 ;
  assign n23714 = n33149 & n23713 ;
  assign n3645 = n2321 & n3639 ;
  assign n2184 = x[107] & n2179 ;
  assign n2258 = x[108] & n2244 ;
  assign n23715 = n2184 | n2258 ;
  assign n23716 = x[109] & n2175 ;
  assign n23717 = n23715 | n23716 ;
  assign n23718 = n3645 | n23717 ;
  assign n33150 = ~n23718 ;
  assign n23719 = x[47] & n33150 ;
  assign n23720 = n29621 & n23718 ;
  assign n23721 = n23719 | n23720 ;
  assign n33151 = ~n23721 ;
  assign n23722 = n23714 & n33151 ;
  assign n33152 = ~n23714 ;
  assign n23723 = n33152 & n23721 ;
  assign n23724 = n23722 | n23723 ;
  assign n33153 = ~n23724 ;
  assign n23725 = n23631 & n33153 ;
  assign n33154 = ~n23631 ;
  assign n23726 = n33154 & n23724 ;
  assign n23727 = n23725 | n23726 ;
  assign n4449 = n2635 & n4442 ;
  assign n2499 = x[110] & n2492 ;
  assign n2566 = x[111] & n2557 ;
  assign n23728 = n2499 | n2566 ;
  assign n23729 = x[112] & n2488 ;
  assign n23730 = n23728 | n23729 ;
  assign n23731 = n4449 | n23730 ;
  assign n33155 = ~n23731 ;
  assign n23732 = x[44] & n33155 ;
  assign n23733 = n29400 & n23731 ;
  assign n23734 = n23732 | n23733 ;
  assign n23735 = n23727 | n23734 ;
  assign n23736 = n23727 & n23734 ;
  assign n33156 = ~n23736 ;
  assign n23737 = n23735 & n33156 ;
  assign n33157 = ~n23547 ;
  assign n23738 = n23456 & n33157 ;
  assign n33158 = ~n23550 ;
  assign n23739 = n33158 & n23557 ;
  assign n23740 = n23738 | n23739 ;
  assign n23741 = n23737 | n23740 ;
  assign n23742 = n23737 & n23740 ;
  assign n33159 = ~n23742 ;
  assign n23743 = n23741 & n33159 ;
  assign n4482 = n3162 & n4474 ;
  assign n3038 = x[113] & n3031 ;
  assign n3108 = x[114] & n3096 ;
  assign n23744 = n3038 | n3108 ;
  assign n23745 = x[115] & n3027 ;
  assign n23746 = n23744 | n23745 ;
  assign n23747 = n4482 | n23746 ;
  assign n33160 = ~n23747 ;
  assign n23748 = x[41] & n33160 ;
  assign n23749 = n29184 & n23747 ;
  assign n23750 = n23748 | n23749 ;
  assign n33161 = ~n23743 ;
  assign n23751 = n33161 & n23750 ;
  assign n33162 = ~n23750 ;
  assign n23752 = n23743 & n33162 ;
  assign n23753 = n23751 | n23752 ;
  assign n23754 = n23629 & n23753 ;
  assign n33163 = ~n23752 ;
  assign n23755 = n23629 & n33163 ;
  assign n23756 = n23751 | n23755 ;
  assign n23757 = n23752 | n23756 ;
  assign n33164 = ~n23754 ;
  assign n23758 = n33164 & n23757 ;
  assign n3594 = n784 & n3574 ;
  assign n3446 = x[116] & n3443 ;
  assign n3538 = x[117] & n3508 ;
  assign n23759 = n3446 | n3538 ;
  assign n23760 = x[118] & n3439 ;
  assign n23761 = n23759 | n23760 ;
  assign n23762 = n3594 | n23761 ;
  assign n33165 = ~n23762 ;
  assign n23763 = x[38] & n33165 ;
  assign n23764 = n28996 & n23762 ;
  assign n23765 = n23763 | n23764 ;
  assign n33166 = ~n23765 ;
  assign n23766 = n23758 & n33166 ;
  assign n33167 = ~n23758 ;
  assign n23767 = n33167 & n23765 ;
  assign n23768 = n23766 | n23767 ;
  assign n23769 = n23627 | n23768 ;
  assign n23770 = n23627 & n23768 ;
  assign n33168 = ~n23770 ;
  assign n23771 = n23769 & n33168 ;
  assign n4986 = n4041 & n4985 ;
  assign n3913 = x[119] & n3910 ;
  assign n3976 = x[120] & n3975 ;
  assign n23772 = n3913 | n3976 ;
  assign n23773 = x[121] & n3906 ;
  assign n23774 = n23772 | n23773 ;
  assign n23775 = n4986 | n23774 ;
  assign n33169 = ~n23775 ;
  assign n23776 = x[35] & n33169 ;
  assign n23777 = n28822 & n23775 ;
  assign n23778 = n23776 | n23777 ;
  assign n23779 = n23771 | n23778 ;
  assign n23780 = n23771 & n23778 ;
  assign n33170 = ~n23780 ;
  assign n23781 = n23779 & n33170 ;
  assign n33171 = ~n23593 ;
  assign n23782 = n23450 & n33171 ;
  assign n23783 = n23592 | n23782 ;
  assign n23784 = n23781 | n23783 ;
  assign n23785 = n23781 & n23783 ;
  assign n33172 = ~n23785 ;
  assign n23786 = n23784 & n33172 ;
  assign n5839 = n779 & n5838 ;
  assign n718 = x[122] & n663 ;
  assign n754 = x[123] & n720 ;
  assign n23787 = n718 | n754 ;
  assign n23788 = x[124] & n652 ;
  assign n23789 = n23787 | n23788 ;
  assign n23790 = n5839 | n23789 ;
  assign n33173 = ~n23790 ;
  assign n23791 = x[32] & n33173 ;
  assign n23792 = n28658 & n23790 ;
  assign n23793 = n23791 | n23792 ;
  assign n23794 = n23438 & n23440 ;
  assign n33174 = ~n23596 ;
  assign n23795 = n23443 & n33174 ;
  assign n23796 = n23794 | n23795 ;
  assign n23797 = n23793 | n23796 ;
  assign n23798 = n23793 & n23796 ;
  assign n33175 = ~n23798 ;
  assign n23799 = n23797 & n33175 ;
  assign n33176 = ~n23786 ;
  assign n23800 = n33176 & n23799 ;
  assign n33177 = ~n23799 ;
  assign n23801 = n23786 & n33177 ;
  assign n23802 = n23800 | n23801 ;
  assign n23803 = n23625 & n23802 ;
  assign n23804 = n23625 | n23802 ;
  assign n33178 = ~n23803 ;
  assign n23805 = n33178 & n23804 ;
  assign n33179 = ~n23805 ;
  assign n23806 = n23613 & n33179 ;
  assign n33180 = ~n23613 ;
  assign n23807 = n33180 & n23805 ;
  assign n23808 = n23806 | n23807 ;
  assign n23809 = n23409 & n23605 ;
  assign n23810 = n23610 | n23809 ;
  assign n23811 = n23808 & n23810 ;
  assign n23812 = n23808 | n23810 ;
  assign n33181 = ~n23811 ;
  assign n219 = n33181 & n23812 ;
  assign n23814 = n23798 | n23800 ;
  assign n6190 = n4632 & n6186 ;
  assign n23815 = x[126] & n4514 ;
  assign n23816 = x[127] & n4572 ;
  assign n23817 = n23815 | n23816 ;
  assign n23818 = n6190 | n23817 ;
  assign n33182 = ~n23818 ;
  assign n23819 = x[29] & n33182 ;
  assign n23820 = n28483 & n23818 ;
  assign n23821 = n23819 | n23820 ;
  assign n23822 = n23814 | n23821 ;
  assign n23823 = n23814 & n23821 ;
  assign n33183 = ~n23823 ;
  assign n23824 = n23822 & n33183 ;
  assign n780 = n642 & n779 ;
  assign n719 = x[123] & n663 ;
  assign n775 = x[124] & n720 ;
  assign n23825 = n719 | n775 ;
  assign n23826 = x[125] & n652 ;
  assign n23827 = n23825 | n23826 ;
  assign n23828 = n780 | n23827 ;
  assign n33184 = ~n23828 ;
  assign n23829 = x[32] & n33184 ;
  assign n23830 = n28658 & n23828 ;
  assign n23831 = n23829 | n23830 ;
  assign n33185 = ~n23771 ;
  assign n23832 = n33185 & n23778 ;
  assign n33186 = ~n23781 ;
  assign n23833 = n33186 & n23783 ;
  assign n23834 = n23832 | n23833 ;
  assign n23835 = n23831 | n23834 ;
  assign n23836 = n23831 & n23834 ;
  assign n33187 = ~n23836 ;
  assign n23837 = n23835 & n33187 ;
  assign n33188 = ~n23768 ;
  assign n23838 = n23627 & n33188 ;
  assign n23839 = n23767 | n23838 ;
  assign n33189 = ~n23685 ;
  assign n23840 = n33189 & n23692 ;
  assign n23841 = n23700 | n23840 ;
  assign n3009 = n1690 & n3001 ;
  assign n1565 = x[102] & n1551 ;
  assign n1632 = x[103] & n1616 ;
  assign n23891 = n1565 | n1632 ;
  assign n23892 = x[104] & n1547 ;
  assign n23893 = n23891 | n23892 ;
  assign n23894 = n3009 | n23893 ;
  assign n23895 = x[53] | n23894 ;
  assign n23896 = x[53] & n23894 ;
  assign n33190 = ~n23896 ;
  assign n23897 = n23895 & n33190 ;
  assign n33191 = ~n23669 ;
  assign n23842 = n33191 & n23676 ;
  assign n23843 = n23684 | n23842 ;
  assign n282 = x[91] & n27215 ;
  assign n853 = x[92] & n805 ;
  assign n23844 = n282 | n853 ;
  assign n23845 = n23649 | n23651 ;
  assign n23846 = n23844 | n23845 ;
  assign n23847 = n23844 & n23845 ;
  assign n33192 = ~n23847 ;
  assign n23848 = n23846 & n33192 ;
  assign n2158 = n1006 & n2152 ;
  assign n907 = x[93] & n900 ;
  assign n980 = x[94] & n949 ;
  assign n23849 = n907 | n980 ;
  assign n23850 = x[95] & n881 ;
  assign n23851 = n23849 | n23850 ;
  assign n23852 = n2158 | n23851 ;
  assign n33193 = ~n23852 ;
  assign n23853 = x[62] & n33193 ;
  assign n23854 = n30886 & n23852 ;
  assign n23855 = n23853 | n23854 ;
  assign n23856 = n23848 | n23855 ;
  assign n23857 = n23848 & n23855 ;
  assign n33194 = ~n23857 ;
  assign n23858 = n23856 & n33194 ;
  assign n33195 = ~n23656 ;
  assign n23859 = n33195 & n23663 ;
  assign n23860 = n23654 | n23859 ;
  assign n23861 = n23858 | n23860 ;
  assign n23862 = n23858 & n23860 ;
  assign n33196 = ~n23862 ;
  assign n23863 = n23861 & n33196 ;
  assign n2849 = n1217 & n2841 ;
  assign n1121 = x[96] & n1079 ;
  assign n1187 = x[97] & n1144 ;
  assign n23864 = n1121 | n1187 ;
  assign n23865 = x[98] & n1075 ;
  assign n23866 = n23864 | n23865 ;
  assign n23867 = n2849 | n23866 ;
  assign n33197 = ~n23867 ;
  assign n23868 = x[59] & n33197 ;
  assign n23869 = n30638 & n23867 ;
  assign n23870 = n23868 | n23869 ;
  assign n23871 = n23863 | n23870 ;
  assign n23872 = n23863 & n23870 ;
  assign n33198 = ~n23872 ;
  assign n23873 = n23871 & n33198 ;
  assign n23874 = n23639 & n23640 ;
  assign n33199 = ~n23666 ;
  assign n23875 = n23643 & n33199 ;
  assign n23876 = n23874 | n23875 ;
  assign n23877 = n23873 | n23876 ;
  assign n23878 = n23873 & n23876 ;
  assign n33200 = ~n23878 ;
  assign n23879 = n23877 & n33200 ;
  assign n2984 = n1457 & n2977 ;
  assign n1341 = x[99] & n1319 ;
  assign n1444 = x[100] & n1384 ;
  assign n23880 = n1341 | n1444 ;
  assign n23881 = x[101] & n1315 ;
  assign n23882 = n23880 | n23881 ;
  assign n23883 = n2984 | n23882 ;
  assign n33201 = ~n23883 ;
  assign n23884 = x[56] & n33201 ;
  assign n23885 = n30379 & n23883 ;
  assign n23886 = n23884 | n23885 ;
  assign n23887 = n23879 | n23886 ;
  assign n23888 = n23879 & n23886 ;
  assign n33202 = ~n23888 ;
  assign n23889 = n23887 & n33202 ;
  assign n23890 = n23843 & n23889 ;
  assign n23898 = n23843 | n23889 ;
  assign n33203 = ~n23890 ;
  assign n23899 = n33203 & n23898 ;
  assign n33204 = ~n23899 ;
  assign n23900 = n23897 & n33204 ;
  assign n33205 = ~n23897 ;
  assign n23901 = n33205 & n23898 ;
  assign n23902 = n33203 & n23901 ;
  assign n23903 = n23900 | n23902 ;
  assign n33206 = ~n23841 ;
  assign n23904 = n33206 & n23903 ;
  assign n33207 = ~n23903 ;
  assign n23905 = n23841 & n33207 ;
  assign n23906 = n23904 | n23905 ;
  assign n3205 = n2007 & n3199 ;
  assign n1885 = x[105] & n1866 ;
  assign n1946 = x[106] & n1931 ;
  assign n23907 = n1885 | n1946 ;
  assign n23908 = x[107] & n1862 ;
  assign n23909 = n23907 | n23908 ;
  assign n23910 = n3205 | n23909 ;
  assign n33208 = ~n23910 ;
  assign n23911 = x[50] & n33208 ;
  assign n23912 = n29865 & n23910 ;
  assign n23913 = n23911 | n23912 ;
  assign n23914 = n23906 | n23913 ;
  assign n23915 = n23906 & n23913 ;
  assign n33209 = ~n23915 ;
  assign n23916 = n23914 & n33209 ;
  assign n33210 = ~n23701 ;
  assign n23917 = n33210 & n23708 ;
  assign n33211 = ~n23711 ;
  assign n23918 = n23632 & n33211 ;
  assign n23919 = n23917 | n23918 ;
  assign n23920 = n23916 | n23919 ;
  assign n23921 = n23916 & n23919 ;
  assign n33212 = ~n23921 ;
  assign n23922 = n23920 & n33212 ;
  assign n3618 = n2321 & n3615 ;
  assign n2187 = x[108] & n2179 ;
  assign n2256 = x[109] & n2244 ;
  assign n23923 = n2187 | n2256 ;
  assign n23924 = x[110] & n2175 ;
  assign n23925 = n23923 | n23924 ;
  assign n23926 = n3618 | n23925 ;
  assign n33213 = ~n23926 ;
  assign n23927 = x[47] & n33213 ;
  assign n23928 = n29621 & n23926 ;
  assign n23929 = n23927 | n23928 ;
  assign n23930 = n23922 | n23929 ;
  assign n23931 = n23922 & n23929 ;
  assign n33214 = ~n23931 ;
  assign n23932 = n23930 & n33214 ;
  assign n23933 = n23723 | n23725 ;
  assign n33215 = ~n23933 ;
  assign n23934 = n23932 & n33215 ;
  assign n33216 = ~n23932 ;
  assign n23935 = n33216 & n23933 ;
  assign n23936 = n23934 | n23935 ;
  assign n4095 = n2635 & n4087 ;
  assign n2498 = x[111] & n2492 ;
  assign n2579 = x[112] & n2557 ;
  assign n23937 = n2498 | n2579 ;
  assign n23938 = x[113] & n2488 ;
  assign n23939 = n23937 | n23938 ;
  assign n23940 = n4095 | n23939 ;
  assign n33217 = ~n23940 ;
  assign n23941 = x[44] & n33217 ;
  assign n23942 = n29400 & n23940 ;
  assign n23943 = n23941 | n23942 ;
  assign n23944 = n23936 | n23943 ;
  assign n23945 = n23936 & n23943 ;
  assign n33218 = ~n23945 ;
  assign n23946 = n23944 & n33218 ;
  assign n33219 = ~n23727 ;
  assign n23947 = n33219 & n23734 ;
  assign n33220 = ~n23737 ;
  assign n23948 = n33220 & n23740 ;
  assign n23949 = n23947 | n23948 ;
  assign n33221 = ~n23949 ;
  assign n23950 = n23946 & n33221 ;
  assign n33222 = ~n23946 ;
  assign n23951 = n33222 & n23949 ;
  assign n23952 = n23950 | n23951 ;
  assign n4707 = n3162 & n4702 ;
  assign n3047 = x[114] & n3031 ;
  assign n3107 = x[115] & n3096 ;
  assign n23953 = n3047 | n3107 ;
  assign n23954 = x[116] & n3027 ;
  assign n23955 = n23953 | n23954 ;
  assign n23956 = n4707 | n23955 ;
  assign n33223 = ~n23956 ;
  assign n23957 = x[41] & n33223 ;
  assign n23958 = n29184 & n23956 ;
  assign n23959 = n23957 | n23958 ;
  assign n23960 = n23952 | n23959 ;
  assign n23961 = n23952 & n23959 ;
  assign n33224 = ~n23961 ;
  assign n23962 = n23960 & n33224 ;
  assign n23963 = n23756 & n23962 ;
  assign n23964 = n23756 | n23962 ;
  assign n33225 = ~n23963 ;
  assign n23965 = n33225 & n23964 ;
  assign n5054 = n3574 & n5047 ;
  assign n3472 = x[117] & n3443 ;
  assign n3515 = x[118] & n3508 ;
  assign n23966 = n3472 | n3515 ;
  assign n23967 = x[119] & n3439 ;
  assign n23968 = n23966 | n23967 ;
  assign n23969 = n5054 | n23968 ;
  assign n33226 = ~n23969 ;
  assign n23970 = x[38] & n33226 ;
  assign n23971 = n28996 & n23969 ;
  assign n23972 = n23970 | n23971 ;
  assign n33227 = ~n23972 ;
  assign n23973 = n23965 & n33227 ;
  assign n33228 = ~n23965 ;
  assign n23974 = n33228 & n23972 ;
  assign n23975 = n23973 | n23974 ;
  assign n33229 = ~n23975 ;
  assign n23976 = n23839 & n33229 ;
  assign n33230 = ~n23839 ;
  assign n23977 = n33230 & n23975 ;
  assign n23978 = n23976 | n23977 ;
  assign n5027 = n4041 & n5022 ;
  assign n3915 = x[120] & n3910 ;
  assign n3977 = x[121] & n3975 ;
  assign n23979 = n3915 | n3977 ;
  assign n23980 = x[122] & n3906 ;
  assign n23981 = n23979 | n23980 ;
  assign n23982 = n5027 | n23981 ;
  assign n33231 = ~n23982 ;
  assign n23983 = x[35] & n33231 ;
  assign n23984 = n28822 & n23982 ;
  assign n23985 = n23983 | n23984 ;
  assign n23986 = n23978 | n23985 ;
  assign n23987 = n23978 & n23985 ;
  assign n33232 = ~n23987 ;
  assign n23988 = n23986 & n33232 ;
  assign n33233 = ~n23988 ;
  assign n23989 = n23837 & n33233 ;
  assign n33234 = ~n23837 ;
  assign n23990 = n33234 & n23988 ;
  assign n33235 = ~n23990 ;
  assign n23991 = n23824 & n33235 ;
  assign n33236 = ~n23989 ;
  assign n23992 = n33236 & n23991 ;
  assign n33237 = ~n23992 ;
  assign n23994 = n23824 & n33237 ;
  assign n23993 = n23990 | n23992 ;
  assign n23995 = n23989 | n23993 ;
  assign n33238 = ~n23994 ;
  assign n23996 = n33238 & n23995 ;
  assign n23997 = n23615 & n23622 ;
  assign n33239 = ~n23802 ;
  assign n23998 = n23625 & n33239 ;
  assign n23999 = n23997 | n23998 ;
  assign n24000 = n23996 | n23999 ;
  assign n24001 = n23996 & n23999 ;
  assign n33240 = ~n24001 ;
  assign n24002 = n24000 & n33240 ;
  assign n24003 = n23613 | n23805 ;
  assign n24004 = n33181 & n24003 ;
  assign n24005 = n24002 & n24004 ;
  assign n24006 = n24002 | n24004 ;
  assign n33241 = ~n24005 ;
  assign n220 = n33241 & n24006 ;
  assign n33242 = ~n23996 ;
  assign n24008 = n33242 & n23999 ;
  assign n33243 = ~n24008 ;
  assign n24009 = n24006 & n33243 ;
  assign n24010 = n23823 | n23992 ;
  assign n24011 = n23836 | n23989 ;
  assign n4571 = x[127] & n4514 ;
  assign n5365 = n4632 & n5360 ;
  assign n24012 = n4571 | n5365 ;
  assign n33244 = ~n24012 ;
  assign n24013 = x[29] & n33244 ;
  assign n24014 = n28483 & n24012 ;
  assign n24015 = n24013 | n24014 ;
  assign n24016 = n24011 | n24015 ;
  assign n24017 = n24011 & n24015 ;
  assign n33245 = ~n24017 ;
  assign n24018 = n24016 & n33245 ;
  assign n5393 = n779 & n5388 ;
  assign n679 = x[124] & n663 ;
  assign n771 = x[125] & n720 ;
  assign n24019 = n679 | n771 ;
  assign n24020 = x[126] & n652 ;
  assign n24021 = n24019 | n24020 ;
  assign n24022 = n5393 | n24021 ;
  assign n33246 = ~n24022 ;
  assign n24023 = x[32] & n33246 ;
  assign n24024 = n28658 & n24022 ;
  assign n24025 = n24023 | n24024 ;
  assign n33247 = ~n23978 ;
  assign n24026 = n33247 & n23985 ;
  assign n24027 = n23976 | n24026 ;
  assign n24028 = n24025 | n24027 ;
  assign n24029 = n24025 & n24027 ;
  assign n33248 = ~n24029 ;
  assign n24030 = n24028 & n33248 ;
  assign n33249 = ~n23962 ;
  assign n24031 = n23756 & n33249 ;
  assign n24032 = n23974 | n24031 ;
  assign n4680 = n3574 & n4678 ;
  assign n3461 = x[118] & n3443 ;
  assign n3512 = x[119] & n3508 ;
  assign n24033 = n3461 | n3512 ;
  assign n24034 = x[120] & n3439 ;
  assign n24035 = n24033 | n24034 ;
  assign n24036 = n4680 | n24035 ;
  assign n33250 = ~n24036 ;
  assign n24037 = x[38] & n33250 ;
  assign n24038 = n28996 & n24036 ;
  assign n24039 = n24037 | n24038 ;
  assign n33251 = ~n23952 ;
  assign n24040 = n33251 & n23959 ;
  assign n24041 = n23951 | n24040 ;
  assign n3193 = n797 & n3162 ;
  assign n3037 = x[115] & n3031 ;
  assign n3105 = x[116] & n3096 ;
  assign n24156 = n3037 | n3105 ;
  assign n24157 = x[117] & n3027 ;
  assign n24158 = n24156 | n24157 ;
  assign n24159 = n3193 | n24158 ;
  assign n24160 = x[41] | n24159 ;
  assign n24161 = x[41] & n24159 ;
  assign n33252 = ~n24161 ;
  assign n24162 = n24160 & n33252 ;
  assign n33253 = ~n23936 ;
  assign n24042 = n33253 & n23943 ;
  assign n24043 = n23935 | n24042 ;
  assign n33254 = ~n23906 ;
  assign n24044 = n33254 & n23913 ;
  assign n24045 = n23905 | n24044 ;
  assign n3882 = n2007 & n3876 ;
  assign n1875 = x[106] & n1866 ;
  assign n1942 = x[107] & n1931 ;
  assign n24046 = n1875 | n1942 ;
  assign n24047 = x[108] & n1862 ;
  assign n24048 = n24046 | n24047 ;
  assign n24049 = n3882 | n24048 ;
  assign n33255 = ~n24049 ;
  assign n24050 = x[50] & n33255 ;
  assign n24051 = n29865 & n24049 ;
  assign n24052 = n24050 | n24051 ;
  assign n33256 = ~n23889 ;
  assign n24053 = n23843 & n33256 ;
  assign n24054 = n23900 | n24053 ;
  assign n33257 = ~n23858 ;
  assign n24055 = n33257 & n23860 ;
  assign n33258 = ~n23863 ;
  assign n24056 = n33258 & n23870 ;
  assign n24057 = n24055 | n24056 ;
  assign n2319 = n1217 & n2313 ;
  assign n1098 = x[97] & n1079 ;
  assign n1164 = x[98] & n1144 ;
  assign n24058 = n1098 | n1164 ;
  assign n24059 = x[99] & n1075 ;
  assign n24060 = n24058 | n24059 ;
  assign n24061 = n2319 | n24060 ;
  assign n33259 = ~n24061 ;
  assign n24062 = x[59] & n33259 ;
  assign n24063 = n30638 & n24061 ;
  assign n24064 = n24062 | n24063 ;
  assign n33260 = ~n23844 ;
  assign n24065 = n33260 & n23845 ;
  assign n33261 = ~n23848 ;
  assign n24066 = n33261 & n23855 ;
  assign n24067 = n24065 | n24066 ;
  assign n283 = x[92] & n27215 ;
  assign n845 = x[93] & n805 ;
  assign n24068 = n283 | n845 ;
  assign n24069 = n33260 & n24068 ;
  assign n33262 = ~n24068 ;
  assign n24070 = n23844 & n33262 ;
  assign n24071 = n24069 | n24070 ;
  assign n24072 = n24067 & n24071 ;
  assign n33263 = ~n24069 ;
  assign n24073 = n24067 & n33263 ;
  assign n24074 = n24070 | n24073 ;
  assign n24075 = n24069 | n24074 ;
  assign n33264 = ~n24072 ;
  assign n24076 = n33264 & n24075 ;
  assign n2006 = n1006 & n2000 ;
  assign n920 = x[94] & n900 ;
  assign n956 = x[95] & n949 ;
  assign n24077 = n920 | n956 ;
  assign n24078 = x[96] & n881 ;
  assign n24079 = n24077 | n24078 ;
  assign n24080 = n2006 | n24079 ;
  assign n33265 = ~n24080 ;
  assign n24081 = x[62] & n33265 ;
  assign n24082 = n30886 & n24080 ;
  assign n24083 = n24081 | n24082 ;
  assign n33266 = ~n24083 ;
  assign n24084 = n24076 & n33266 ;
  assign n33267 = ~n24076 ;
  assign n24085 = n33267 & n24083 ;
  assign n24086 = n24084 | n24085 ;
  assign n33268 = ~n24064 ;
  assign n24087 = n33268 & n24086 ;
  assign n33269 = ~n24086 ;
  assign n24088 = n24064 & n33269 ;
  assign n24089 = n24087 | n24088 ;
  assign n33270 = ~n24089 ;
  assign n24090 = n24057 & n33270 ;
  assign n33271 = ~n24057 ;
  assign n24091 = n33271 & n24089 ;
  assign n24092 = n24090 | n24091 ;
  assign n2874 = n1457 & n2867 ;
  assign n1354 = x[100] & n1319 ;
  assign n1440 = x[101] & n1384 ;
  assign n24093 = n1354 | n1440 ;
  assign n24094 = x[102] & n1315 ;
  assign n24095 = n24093 | n24094 ;
  assign n24096 = n2874 | n24095 ;
  assign n33272 = ~n24096 ;
  assign n24097 = x[56] & n33272 ;
  assign n24098 = n30379 & n24096 ;
  assign n24099 = n24097 | n24098 ;
  assign n24100 = n24092 | n24099 ;
  assign n24101 = n24092 & n24099 ;
  assign n33273 = ~n24101 ;
  assign n24102 = n24100 & n33273 ;
  assign n33274 = ~n23873 ;
  assign n24103 = n33274 & n23876 ;
  assign n33275 = ~n23879 ;
  assign n24104 = n33275 & n23886 ;
  assign n24105 = n24103 | n24104 ;
  assign n33276 = ~n24105 ;
  assign n24106 = n24102 & n33276 ;
  assign n33277 = ~n24102 ;
  assign n24107 = n33277 & n24105 ;
  assign n24108 = n24106 | n24107 ;
  assign n3418 = n1690 & n3409 ;
  assign n1564 = x[103] & n1551 ;
  assign n1666 = x[104] & n1616 ;
  assign n24109 = n1564 | n1666 ;
  assign n24110 = x[105] & n1547 ;
  assign n24111 = n24109 | n24110 ;
  assign n24112 = n3418 | n24111 ;
  assign n33278 = ~n24112 ;
  assign n24113 = x[53] & n33278 ;
  assign n24114 = n30125 & n24112 ;
  assign n24115 = n24113 | n24114 ;
  assign n33279 = ~n24115 ;
  assign n24116 = n24108 & n33279 ;
  assign n33280 = ~n24108 ;
  assign n24117 = n33280 & n24115 ;
  assign n24118 = n24116 | n24117 ;
  assign n33281 = ~n24054 ;
  assign n24119 = n33281 & n24118 ;
  assign n33282 = ~n24118 ;
  assign n24120 = n24054 & n33282 ;
  assign n24121 = n24119 | n24120 ;
  assign n24122 = n24052 | n24121 ;
  assign n24123 = n24052 & n24121 ;
  assign n33283 = ~n24123 ;
  assign n24124 = n24122 & n33283 ;
  assign n24125 = n24045 | n24124 ;
  assign n24126 = n24045 & n24124 ;
  assign n33284 = ~n24126 ;
  assign n24127 = n24125 & n33284 ;
  assign n4252 = n2321 & n4246 ;
  assign n2183 = x[109] & n2179 ;
  assign n2257 = x[110] & n2244 ;
  assign n24128 = n2183 | n2257 ;
  assign n24129 = x[111] & n2175 ;
  assign n24130 = n24128 | n24129 ;
  assign n24131 = n4252 | n24130 ;
  assign n33285 = ~n24131 ;
  assign n24132 = x[47] & n33285 ;
  assign n24133 = n29621 & n24131 ;
  assign n24134 = n24132 | n24133 ;
  assign n24135 = n24127 | n24134 ;
  assign n24136 = n24127 & n24134 ;
  assign n33286 = ~n24136 ;
  assign n24137 = n24135 & n33286 ;
  assign n33287 = ~n23916 ;
  assign n24138 = n33287 & n23919 ;
  assign n33288 = ~n23922 ;
  assign n24139 = n33288 & n23929 ;
  assign n24140 = n24138 | n24139 ;
  assign n33289 = ~n24140 ;
  assign n24141 = n24137 & n33289 ;
  assign n33290 = ~n24137 ;
  assign n24142 = n33290 & n24140 ;
  assign n24143 = n24141 | n24142 ;
  assign n4283 = n2635 & n4276 ;
  assign n2497 = x[112] & n2492 ;
  assign n2572 = x[113] & n2557 ;
  assign n24144 = n2497 | n2572 ;
  assign n24145 = x[114] & n2488 ;
  assign n24146 = n24144 | n24145 ;
  assign n24147 = n4283 | n24146 ;
  assign n33291 = ~n24147 ;
  assign n24148 = x[44] & n33291 ;
  assign n24149 = n29400 & n24147 ;
  assign n24150 = n24148 | n24149 ;
  assign n24151 = n24143 | n24150 ;
  assign n24152 = n24143 & n24150 ;
  assign n33292 = ~n24152 ;
  assign n24153 = n24151 & n33292 ;
  assign n24154 = n24043 | n24153 ;
  assign n24155 = n24043 & n24153 ;
  assign n33293 = ~n24155 ;
  assign n24163 = n24154 & n33293 ;
  assign n33294 = ~n24163 ;
  assign n24164 = n24162 & n33294 ;
  assign n33295 = ~n24162 ;
  assign n24165 = n24154 & n33295 ;
  assign n24166 = n33293 & n24165 ;
  assign n24167 = n24164 | n24166 ;
  assign n33296 = ~n24041 ;
  assign n24168 = n33296 & n24167 ;
  assign n33297 = ~n24167 ;
  assign n24169 = n24041 & n33297 ;
  assign n24170 = n24168 | n24169 ;
  assign n24171 = n24039 | n24170 ;
  assign n24172 = n24039 & n24170 ;
  assign n33298 = ~n24172 ;
  assign n24173 = n24171 & n33298 ;
  assign n33299 = ~n24173 ;
  assign n24174 = n24032 & n33299 ;
  assign n33300 = ~n24032 ;
  assign n24175 = n33300 & n24173 ;
  assign n24176 = n24174 | n24175 ;
  assign n5419 = n4041 & n5417 ;
  assign n3912 = x[121] & n3910 ;
  assign n4010 = x[122] & n3975 ;
  assign n24177 = n3912 | n4010 ;
  assign n24178 = x[123] & n3906 ;
  assign n24179 = n24177 | n24178 ;
  assign n24180 = n5419 | n24179 ;
  assign n33301 = ~n24180 ;
  assign n24181 = x[35] & n33301 ;
  assign n24182 = n28822 & n24180 ;
  assign n24183 = n24181 | n24182 ;
  assign n24184 = n24176 | n24183 ;
  assign n24185 = n24176 & n24183 ;
  assign n33302 = ~n24185 ;
  assign n24186 = n24184 & n33302 ;
  assign n24187 = n24030 & n24186 ;
  assign n24188 = n24030 | n24186 ;
  assign n33303 = ~n24187 ;
  assign n24189 = n33303 & n24188 ;
  assign n24190 = n24018 | n24189 ;
  assign n24191 = n24018 & n24189 ;
  assign n33304 = ~n24191 ;
  assign n24192 = n24190 & n33304 ;
  assign n24193 = n24010 & n24192 ;
  assign n24194 = n24010 | n24192 ;
  assign n33305 = ~n24193 ;
  assign n24195 = n33305 & n24194 ;
  assign n24196 = n24009 | n24195 ;
  assign n24197 = n24009 & n24194 ;
  assign n24198 = n33305 & n24197 ;
  assign n33306 = ~n24198 ;
  assign n221 = n24196 & n33306 ;
  assign n33307 = ~n24192 ;
  assign n24200 = n24010 & n33307 ;
  assign n33308 = ~n24200 ;
  assign n24201 = n24196 & n33308 ;
  assign n33309 = ~n24189 ;
  assign n24202 = n24018 & n33309 ;
  assign n24203 = n24017 | n24202 ;
  assign n33310 = ~n24153 ;
  assign n24204 = n24043 & n33310 ;
  assign n24205 = n24164 | n24204 ;
  assign n33311 = ~n24143 ;
  assign n24206 = n33311 & n24150 ;
  assign n24207 = n24142 | n24206 ;
  assign n33312 = ~n24121 ;
  assign n24208 = n24052 & n33312 ;
  assign n24209 = n24120 | n24208 ;
  assign n24210 = n24107 | n24117 ;
  assign n24211 = n24085 | n24088 ;
  assign n284 = x[93] & n27215 ;
  assign n860 = x[94] & n805 ;
  assign n24212 = n284 | n860 ;
  assign n33313 = ~n24212 ;
  assign n24213 = x[29] & n33313 ;
  assign n24214 = n28483 & n24212 ;
  assign n24215 = n24213 | n24214 ;
  assign n24216 = n24068 | n24215 ;
  assign n24218 = n24068 & n24215 ;
  assign n33314 = ~n24218 ;
  assign n24219 = n24216 & n33314 ;
  assign n24220 = n24074 & n24219 ;
  assign n24221 = n24074 | n24219 ;
  assign n33315 = ~n24220 ;
  assign n24222 = n33315 & n24221 ;
  assign n2442 = n1006 & n2438 ;
  assign n906 = x[95] & n900 ;
  assign n958 = x[96] & n949 ;
  assign n24223 = n906 | n958 ;
  assign n24224 = x[97] & n881 ;
  assign n24225 = n24223 | n24224 ;
  assign n24226 = n2442 | n24225 ;
  assign n33316 = ~n24226 ;
  assign n24227 = x[62] & n33316 ;
  assign n24228 = n30886 & n24226 ;
  assign n24229 = n24227 | n24228 ;
  assign n33317 = ~n24229 ;
  assign n24230 = n24222 & n33317 ;
  assign n33318 = ~n24222 ;
  assign n24231 = n33318 & n24229 ;
  assign n24232 = n24230 | n24231 ;
  assign n2472 = n1217 & n2466 ;
  assign n1097 = x[98] & n1079 ;
  assign n1163 = x[99] & n1144 ;
  assign n24233 = n1097 | n1163 ;
  assign n24234 = x[100] & n1075 ;
  assign n24235 = n24233 | n24234 ;
  assign n24236 = n2472 | n24235 ;
  assign n33319 = ~n24236 ;
  assign n24237 = x[59] & n33319 ;
  assign n24238 = n30638 & n24236 ;
  assign n24239 = n24237 | n24238 ;
  assign n33320 = ~n24239 ;
  assign n24240 = n24232 & n33320 ;
  assign n33321 = ~n24232 ;
  assign n24241 = n33321 & n24239 ;
  assign n24242 = n24240 | n24241 ;
  assign n33322 = ~n24242 ;
  assign n24243 = n24211 & n33322 ;
  assign n33323 = ~n24211 ;
  assign n24244 = n33323 & n24242 ;
  assign n24245 = n24243 | n24244 ;
  assign n2632 = n1457 & n2626 ;
  assign n1340 = x[101] & n1319 ;
  assign n1404 = x[102] & n1384 ;
  assign n24246 = n1340 | n1404 ;
  assign n24247 = x[103] & n1315 ;
  assign n24248 = n24246 | n24247 ;
  assign n24249 = n2632 | n24248 ;
  assign n33324 = ~n24249 ;
  assign n24250 = x[56] & n33324 ;
  assign n24251 = n30379 & n24249 ;
  assign n24252 = n24250 | n24251 ;
  assign n24253 = n24245 | n24252 ;
  assign n24254 = n24245 & n24252 ;
  assign n33325 = ~n24254 ;
  assign n24255 = n24253 & n33325 ;
  assign n33326 = ~n24092 ;
  assign n24256 = n33326 & n24099 ;
  assign n24257 = n24090 | n24256 ;
  assign n33327 = ~n24257 ;
  assign n24258 = n24255 & n33327 ;
  assign n33328 = ~n24255 ;
  assign n24259 = n33328 & n24257 ;
  assign n24260 = n24258 | n24259 ;
  assign n3226 = n1690 & n3223 ;
  assign n1562 = x[104] & n1551 ;
  assign n1652 = x[105] & n1616 ;
  assign n24261 = n1562 | n1652 ;
  assign n24262 = x[106] & n1547 ;
  assign n24263 = n24261 | n24262 ;
  assign n24264 = n3226 | n24263 ;
  assign n33329 = ~n24264 ;
  assign n24265 = x[53] & n33329 ;
  assign n24266 = n30125 & n24264 ;
  assign n24267 = n24265 | n24266 ;
  assign n24268 = n24260 | n24267 ;
  assign n24269 = n24260 & n24267 ;
  assign n33330 = ~n24269 ;
  assign n24270 = n24268 & n33330 ;
  assign n24271 = n24210 & n24270 ;
  assign n24272 = n24210 | n24270 ;
  assign n33331 = ~n24271 ;
  assign n24273 = n33331 & n24272 ;
  assign n3647 = n2007 & n3639 ;
  assign n1916 = x[107] & n1866 ;
  assign n1944 = x[108] & n1931 ;
  assign n24274 = n1916 | n1944 ;
  assign n24275 = x[109] & n1862 ;
  assign n24276 = n24274 | n24275 ;
  assign n24277 = n3647 | n24276 ;
  assign n33332 = ~n24277 ;
  assign n24278 = x[50] & n33332 ;
  assign n24279 = n29865 & n24277 ;
  assign n24280 = n24278 | n24279 ;
  assign n33333 = ~n24280 ;
  assign n24281 = n24273 & n33333 ;
  assign n33334 = ~n24273 ;
  assign n24282 = n33334 & n24280 ;
  assign n24283 = n24281 | n24282 ;
  assign n33335 = ~n24283 ;
  assign n24284 = n24209 & n33335 ;
  assign n33336 = ~n24209 ;
  assign n24285 = n33336 & n24283 ;
  assign n24286 = n24284 | n24285 ;
  assign n4448 = n2321 & n4442 ;
  assign n2207 = x[110] & n2179 ;
  assign n2283 = x[111] & n2244 ;
  assign n24287 = n2207 | n2283 ;
  assign n24288 = x[112] & n2175 ;
  assign n24289 = n24287 | n24288 ;
  assign n24290 = n4448 | n24289 ;
  assign n33337 = ~n24290 ;
  assign n24291 = x[47] & n33337 ;
  assign n24292 = n29621 & n24290 ;
  assign n24293 = n24291 | n24292 ;
  assign n24294 = n24286 | n24293 ;
  assign n24295 = n24286 & n24293 ;
  assign n33338 = ~n24295 ;
  assign n24296 = n24294 & n33338 ;
  assign n33339 = ~n24124 ;
  assign n24297 = n24045 & n33339 ;
  assign n33340 = ~n24127 ;
  assign n24298 = n33340 & n24134 ;
  assign n24299 = n24297 | n24298 ;
  assign n24300 = n24296 | n24299 ;
  assign n24301 = n24296 & n24299 ;
  assign n33341 = ~n24301 ;
  assign n24302 = n24300 & n33341 ;
  assign n4477 = n2635 & n4474 ;
  assign n2513 = x[113] & n2492 ;
  assign n2563 = x[114] & n2557 ;
  assign n24303 = n2513 | n2563 ;
  assign n24304 = x[115] & n2488 ;
  assign n24305 = n24303 | n24304 ;
  assign n24306 = n4477 | n24305 ;
  assign n33342 = ~n24306 ;
  assign n24307 = x[44] & n33342 ;
  assign n24308 = n29400 & n24306 ;
  assign n24309 = n24307 | n24308 ;
  assign n33343 = ~n24302 ;
  assign n24310 = n33343 & n24309 ;
  assign n33344 = ~n24309 ;
  assign n24311 = n24302 & n33344 ;
  assign n24312 = n24310 | n24311 ;
  assign n24313 = n24207 & n24312 ;
  assign n33345 = ~n24311 ;
  assign n24314 = n24207 & n33345 ;
  assign n24315 = n24310 | n24314 ;
  assign n24316 = n24311 | n24315 ;
  assign n33346 = ~n24313 ;
  assign n24317 = n33346 & n24316 ;
  assign n3164 = n784 & n3162 ;
  assign n3044 = x[116] & n3031 ;
  assign n3148 = x[117] & n3096 ;
  assign n24318 = n3044 | n3148 ;
  assign n24319 = x[118] & n3027 ;
  assign n24320 = n24318 | n24319 ;
  assign n24321 = n3164 | n24320 ;
  assign n33347 = ~n24321 ;
  assign n24322 = x[41] & n33347 ;
  assign n24323 = n29184 & n24321 ;
  assign n24324 = n24322 | n24323 ;
  assign n33348 = ~n24324 ;
  assign n24325 = n24317 & n33348 ;
  assign n33349 = ~n24317 ;
  assign n24326 = n33349 & n24324 ;
  assign n24327 = n24325 | n24326 ;
  assign n24328 = n24205 | n24327 ;
  assign n24329 = n24205 & n24327 ;
  assign n33350 = ~n24329 ;
  assign n24330 = n24328 & n33350 ;
  assign n4988 = n3574 & n4985 ;
  assign n3470 = x[119] & n3443 ;
  assign n3562 = x[120] & n3508 ;
  assign n24331 = n3470 | n3562 ;
  assign n24332 = x[121] & n3439 ;
  assign n24333 = n24331 | n24332 ;
  assign n24334 = n4988 | n24333 ;
  assign n33351 = ~n24334 ;
  assign n24335 = x[38] & n33351 ;
  assign n24336 = n28996 & n24334 ;
  assign n24337 = n24335 | n24336 ;
  assign n24338 = n24330 | n24337 ;
  assign n24339 = n24330 & n24337 ;
  assign n33352 = ~n24339 ;
  assign n24340 = n24338 & n33352 ;
  assign n33353 = ~n24170 ;
  assign n24341 = n24039 & n33353 ;
  assign n24342 = n24169 | n24341 ;
  assign n24343 = n24340 | n24342 ;
  assign n24344 = n24340 & n24342 ;
  assign n33354 = ~n24344 ;
  assign n24345 = n24343 & n33354 ;
  assign n5844 = n4041 & n5838 ;
  assign n3911 = x[122] & n3910 ;
  assign n4021 = x[123] & n3975 ;
  assign n24346 = n3911 | n4021 ;
  assign n24347 = x[124] & n3906 ;
  assign n24348 = n24346 | n24347 ;
  assign n24349 = n5844 | n24348 ;
  assign n33355 = ~n24349 ;
  assign n24350 = x[35] & n33355 ;
  assign n24351 = n28822 & n24349 ;
  assign n24352 = n24350 | n24351 ;
  assign n24353 = n24345 | n24352 ;
  assign n24354 = n24345 & n24352 ;
  assign n33356 = ~n24354 ;
  assign n24355 = n24353 & n33356 ;
  assign n33357 = ~n24176 ;
  assign n24356 = n33357 & n24183 ;
  assign n24357 = n24174 | n24356 ;
  assign n33358 = ~n24357 ;
  assign n24358 = n24355 & n33358 ;
  assign n33359 = ~n24355 ;
  assign n24359 = n33359 & n24357 ;
  assign n24360 = n24358 | n24359 ;
  assign n33360 = ~n24186 ;
  assign n24361 = n24030 & n33360 ;
  assign n24362 = n24029 | n24361 ;
  assign n5631 = n779 & n5629 ;
  assign n669 = x[125] & n663 ;
  assign n758 = x[126] & n720 ;
  assign n24363 = n669 | n758 ;
  assign n24364 = x[127] & n652 ;
  assign n24365 = n24363 | n24364 ;
  assign n24366 = n5631 | n24365 ;
  assign n33361 = ~n24366 ;
  assign n24367 = x[32] & n33361 ;
  assign n24368 = n28658 & n24366 ;
  assign n24369 = n24367 | n24368 ;
  assign n33362 = ~n24369 ;
  assign n24370 = n24362 & n33362 ;
  assign n33363 = ~n24362 ;
  assign n24371 = n33363 & n24369 ;
  assign n24372 = n24370 | n24371 ;
  assign n24373 = n24360 | n24372 ;
  assign n24374 = n24360 & n24372 ;
  assign n33364 = ~n24374 ;
  assign n24375 = n24373 & n33364 ;
  assign n24376 = n24203 | n24375 ;
  assign n24377 = n24203 & n24375 ;
  assign n33365 = ~n24377 ;
  assign n24378 = n24376 & n33365 ;
  assign n24379 = n24201 & n24378 ;
  assign n24380 = n24201 | n24378 ;
  assign n33366 = ~n24379 ;
  assign n222 = n33366 & n24380 ;
  assign n33367 = ~n24345 ;
  assign n24532 = n33367 & n24352 ;
  assign n24533 = n24359 | n24532 ;
  assign n6192 = n779 & n6186 ;
  assign n24534 = x[126] & n663 ;
  assign n24535 = x[127] & n720 ;
  assign n24536 = n24534 | n24535 ;
  assign n24537 = n6192 | n24536 ;
  assign n33368 = ~n24537 ;
  assign n24538 = x[32] & n33368 ;
  assign n24539 = n28658 & n24537 ;
  assign n24540 = n24538 | n24539 ;
  assign n24541 = n24533 | n24540 ;
  assign n24542 = n24533 & n24540 ;
  assign n33369 = ~n24542 ;
  assign n24543 = n24541 & n33369 ;
  assign n33370 = ~n24327 ;
  assign n24382 = n24205 & n33370 ;
  assign n24383 = n24326 | n24382 ;
  assign n33371 = ~n24245 ;
  assign n24384 = n33371 & n24252 ;
  assign n24385 = n24259 | n24384 ;
  assign n3010 = n1457 & n3001 ;
  assign n1325 = x[102] & n1319 ;
  assign n1409 = x[103] & n1384 ;
  assign n24420 = n1325 | n1409 ;
  assign n24421 = x[104] & n1315 ;
  assign n24422 = n24420 | n24421 ;
  assign n24423 = n3010 | n24422 ;
  assign n24424 = x[56] | n24423 ;
  assign n24425 = x[56] & n24423 ;
  assign n33372 = ~n24425 ;
  assign n24426 = n24424 & n33372 ;
  assign n24386 = n24241 | n24243 ;
  assign n2985 = n1217 & n2977 ;
  assign n1124 = x[99] & n1079 ;
  assign n1161 = x[100] & n1144 ;
  assign n24406 = n1124 | n1161 ;
  assign n24407 = x[101] & n1075 ;
  assign n24408 = n24406 | n24407 ;
  assign n24409 = n2985 | n24408 ;
  assign n24410 = x[59] | n24409 ;
  assign n24411 = x[59] & n24409 ;
  assign n33373 = ~n24411 ;
  assign n24412 = n24410 & n33373 ;
  assign n33374 = ~n24219 ;
  assign n24387 = n24074 & n33374 ;
  assign n24388 = n24231 | n24387 ;
  assign n285 = x[94] & n27215 ;
  assign n840 = x[95] & n805 ;
  assign n24389 = n285 | n840 ;
  assign n33375 = ~n24215 ;
  assign n24217 = n24068 & n33375 ;
  assign n24390 = n24214 | n24217 ;
  assign n24391 = n24389 | n24390 ;
  assign n24392 = n24389 & n24390 ;
  assign n33376 = ~n24392 ;
  assign n24393 = n24391 & n33376 ;
  assign n2850 = n1006 & n2841 ;
  assign n905 = x[96] & n900 ;
  assign n955 = x[97] & n949 ;
  assign n24394 = n905 | n955 ;
  assign n24395 = x[98] & n881 ;
  assign n24396 = n24394 | n24395 ;
  assign n24397 = n2850 | n24396 ;
  assign n33377 = ~n24397 ;
  assign n24398 = x[62] & n33377 ;
  assign n24399 = n30886 & n24397 ;
  assign n24400 = n24398 | n24399 ;
  assign n24401 = n24393 | n24400 ;
  assign n24402 = n24393 & n24400 ;
  assign n33378 = ~n24402 ;
  assign n24403 = n24401 & n33378 ;
  assign n24405 = n24388 & n24403 ;
  assign n24413 = n24388 | n24403 ;
  assign n33379 = ~n24405 ;
  assign n24414 = n33379 & n24413 ;
  assign n33380 = ~n24414 ;
  assign n24415 = n24412 & n33380 ;
  assign n33381 = ~n24412 ;
  assign n24416 = n33381 & n24413 ;
  assign n24417 = n33379 & n24416 ;
  assign n24418 = n24415 | n24417 ;
  assign n24419 = n24386 & n24418 ;
  assign n24427 = n24386 | n24418 ;
  assign n33382 = ~n24419 ;
  assign n24428 = n33382 & n24427 ;
  assign n33383 = ~n24428 ;
  assign n24429 = n24426 & n33383 ;
  assign n33384 = ~n24426 ;
  assign n24430 = n33384 & n24427 ;
  assign n24431 = n33382 & n24430 ;
  assign n24432 = n24429 | n24431 ;
  assign n33385 = ~n24385 ;
  assign n24433 = n33385 & n24432 ;
  assign n33386 = ~n24432 ;
  assign n24434 = n24385 & n33386 ;
  assign n24435 = n24433 | n24434 ;
  assign n3207 = n1690 & n3199 ;
  assign n1561 = x[105] & n1551 ;
  assign n1631 = x[106] & n1616 ;
  assign n24436 = n1561 | n1631 ;
  assign n24437 = x[107] & n1547 ;
  assign n24438 = n24436 | n24437 ;
  assign n24439 = n3207 | n24438 ;
  assign n33387 = ~n24439 ;
  assign n24440 = x[53] & n33387 ;
  assign n24441 = n30125 & n24439 ;
  assign n24442 = n24440 | n24441 ;
  assign n24443 = n24435 | n24442 ;
  assign n24444 = n24435 & n24442 ;
  assign n33388 = ~n24444 ;
  assign n24445 = n24443 & n33388 ;
  assign n33389 = ~n24260 ;
  assign n24446 = n33389 & n24267 ;
  assign n33390 = ~n24270 ;
  assign n24447 = n24210 & n33390 ;
  assign n24448 = n24446 | n24447 ;
  assign n24449 = n24445 | n24448 ;
  assign n24450 = n24445 & n24448 ;
  assign n33391 = ~n24450 ;
  assign n24451 = n24449 & n33391 ;
  assign n3620 = n2007 & n3615 ;
  assign n1924 = x[108] & n1866 ;
  assign n1941 = x[109] & n1931 ;
  assign n24452 = n1924 | n1941 ;
  assign n24453 = x[110] & n1862 ;
  assign n24454 = n24452 | n24453 ;
  assign n24455 = n3620 | n24454 ;
  assign n33392 = ~n24455 ;
  assign n24456 = x[50] & n33392 ;
  assign n24457 = n29865 & n24455 ;
  assign n24458 = n24456 | n24457 ;
  assign n24459 = n24451 | n24458 ;
  assign n24460 = n24451 & n24458 ;
  assign n33393 = ~n24460 ;
  assign n24461 = n24459 & n33393 ;
  assign n24462 = n24282 | n24284 ;
  assign n33394 = ~n24462 ;
  assign n24463 = n24461 & n33394 ;
  assign n33395 = ~n24461 ;
  assign n24464 = n33395 & n24462 ;
  assign n24465 = n24463 | n24464 ;
  assign n4093 = n2321 & n4087 ;
  assign n2196 = x[111] & n2179 ;
  assign n2255 = x[112] & n2244 ;
  assign n24466 = n2196 | n2255 ;
  assign n24467 = x[113] & n2175 ;
  assign n24468 = n24466 | n24467 ;
  assign n24469 = n4093 | n24468 ;
  assign n33396 = ~n24469 ;
  assign n24470 = x[47] & n33396 ;
  assign n24471 = n29621 & n24469 ;
  assign n24472 = n24470 | n24471 ;
  assign n24473 = n24465 | n24472 ;
  assign n24474 = n24465 & n24472 ;
  assign n33397 = ~n24474 ;
  assign n24475 = n24473 & n33397 ;
  assign n33398 = ~n24286 ;
  assign n24476 = n33398 & n24293 ;
  assign n33399 = ~n24296 ;
  assign n24477 = n33399 & n24299 ;
  assign n24478 = n24476 | n24477 ;
  assign n33400 = ~n24478 ;
  assign n24479 = n24475 & n33400 ;
  assign n33401 = ~n24475 ;
  assign n24480 = n33401 & n24478 ;
  assign n24481 = n24479 | n24480 ;
  assign n4709 = n2635 & n4702 ;
  assign n2495 = x[114] & n2492 ;
  assign n2561 = x[115] & n2557 ;
  assign n24482 = n2495 | n2561 ;
  assign n24483 = x[116] & n2488 ;
  assign n24484 = n24482 | n24483 ;
  assign n24485 = n4709 | n24484 ;
  assign n33402 = ~n24485 ;
  assign n24486 = x[44] & n33402 ;
  assign n24487 = n29400 & n24485 ;
  assign n24488 = n24486 | n24487 ;
  assign n24489 = n24481 | n24488 ;
  assign n24490 = n24481 & n24488 ;
  assign n33403 = ~n24490 ;
  assign n24491 = n24489 & n33403 ;
  assign n24492 = n24315 & n24491 ;
  assign n24493 = n24315 | n24491 ;
  assign n33404 = ~n24492 ;
  assign n24494 = n33404 & n24493 ;
  assign n5051 = n3162 & n5047 ;
  assign n3035 = x[117] & n3031 ;
  assign n3102 = x[118] & n3096 ;
  assign n24495 = n3035 | n3102 ;
  assign n24496 = x[119] & n3027 ;
  assign n24497 = n24495 | n24496 ;
  assign n24498 = n5051 | n24497 ;
  assign n33405 = ~n24498 ;
  assign n24499 = x[41] & n33405 ;
  assign n24500 = n29184 & n24498 ;
  assign n24501 = n24499 | n24500 ;
  assign n33406 = ~n24501 ;
  assign n24502 = n24494 & n33406 ;
  assign n33407 = ~n24494 ;
  assign n24503 = n33407 & n24501 ;
  assign n24504 = n24502 | n24503 ;
  assign n33408 = ~n24504 ;
  assign n24505 = n24383 & n33408 ;
  assign n33409 = ~n24383 ;
  assign n24506 = n33409 & n24504 ;
  assign n24507 = n24505 | n24506 ;
  assign n5026 = n3574 & n5022 ;
  assign n3481 = x[120] & n3443 ;
  assign n3509 = x[121] & n3508 ;
  assign n24508 = n3481 | n3509 ;
  assign n24509 = x[122] & n3439 ;
  assign n24510 = n24508 | n24509 ;
  assign n24511 = n5026 | n24510 ;
  assign n33410 = ~n24511 ;
  assign n24512 = x[38] & n33410 ;
  assign n24513 = n28996 & n24511 ;
  assign n24514 = n24512 | n24513 ;
  assign n24515 = n24507 | n24514 ;
  assign n24516 = n24507 & n24514 ;
  assign n33411 = ~n24516 ;
  assign n24517 = n24515 & n33411 ;
  assign n33412 = ~n24330 ;
  assign n24518 = n33412 & n24337 ;
  assign n33413 = ~n24340 ;
  assign n24519 = n33413 & n24342 ;
  assign n24520 = n24518 | n24519 ;
  assign n33414 = ~n24520 ;
  assign n24521 = n24517 & n33414 ;
  assign n33415 = ~n24517 ;
  assign n24522 = n33415 & n24520 ;
  assign n24523 = n24521 | n24522 ;
  assign n4083 = n642 & n4041 ;
  assign n3970 = x[123] & n3910 ;
  assign n4037 = x[124] & n3975 ;
  assign n24524 = n3970 | n4037 ;
  assign n24525 = x[125] & n3906 ;
  assign n24526 = n24524 | n24525 ;
  assign n24527 = n4083 | n24526 ;
  assign n33416 = ~n24527 ;
  assign n24528 = x[35] & n33416 ;
  assign n24529 = n28822 & n24527 ;
  assign n24530 = n24528 | n24529 ;
  assign n33417 = ~n24523 ;
  assign n24531 = n33417 & n24530 ;
  assign n33418 = ~n24530 ;
  assign n24544 = n24523 & n33418 ;
  assign n33419 = ~n24544 ;
  assign n24545 = n24543 & n33419 ;
  assign n33420 = ~n24531 ;
  assign n24546 = n33420 & n24545 ;
  assign n33421 = ~n24546 ;
  assign n24547 = n24543 & n33421 ;
  assign n24548 = n24544 | n24546 ;
  assign n24549 = n24531 | n24548 ;
  assign n33422 = ~n24547 ;
  assign n24550 = n33422 & n24549 ;
  assign n24551 = n24362 & n24369 ;
  assign n33423 = ~n24360 ;
  assign n24552 = n33423 & n24372 ;
  assign n24553 = n24551 | n24552 ;
  assign n33424 = ~n24553 ;
  assign n24554 = n24550 & n33424 ;
  assign n33425 = ~n24550 ;
  assign n24555 = n33425 & n24553 ;
  assign n24556 = n24554 | n24555 ;
  assign n33426 = ~n24375 ;
  assign n24557 = n24203 & n33426 ;
  assign n33427 = ~n24557 ;
  assign n24558 = n24380 & n33427 ;
  assign n24559 = n24556 | n24558 ;
  assign n24560 = n24556 & n24558 ;
  assign n33428 = ~n24560 ;
  assign n223 = n24559 & n33428 ;
  assign n33429 = ~n24555 ;
  assign n24729 = n33429 & n24559 ;
  assign n24562 = n24542 | n24546 ;
  assign n24563 = n24522 | n24531 ;
  assign n716 = x[127] & n663 ;
  assign n5363 = n779 & n5360 ;
  assign n24564 = n716 | n5363 ;
  assign n33430 = ~n24564 ;
  assign n24565 = x[32] & n33430 ;
  assign n24566 = n28658 & n24564 ;
  assign n24567 = n24565 | n24566 ;
  assign n24568 = n24563 | n24567 ;
  assign n24569 = n24563 & n24567 ;
  assign n33431 = ~n24569 ;
  assign n24570 = n24568 & n33431 ;
  assign n33432 = ~n24491 ;
  assign n24571 = n24315 & n33432 ;
  assign n24572 = n24503 | n24571 ;
  assign n4686 = n3162 & n4678 ;
  assign n3084 = x[118] & n3031 ;
  assign n3100 = x[119] & n3096 ;
  assign n24573 = n3084 | n3100 ;
  assign n24574 = x[120] & n3027 ;
  assign n24575 = n24573 | n24574 ;
  assign n24576 = n4686 | n24575 ;
  assign n33433 = ~n24576 ;
  assign n24577 = x[41] & n33433 ;
  assign n24578 = n29184 & n24576 ;
  assign n24579 = n24577 | n24578 ;
  assign n33434 = ~n24481 ;
  assign n24580 = n33434 & n24488 ;
  assign n24581 = n24480 | n24580 ;
  assign n2636 = n797 & n2635 ;
  assign n2532 = x[115] & n2492 ;
  assign n2613 = x[116] & n2557 ;
  assign n24679 = n2532 | n2613 ;
  assign n24680 = x[117] & n2488 ;
  assign n24681 = n24679 | n24680 ;
  assign n24682 = n2636 | n24681 ;
  assign n24683 = x[44] | n24682 ;
  assign n24684 = x[44] & n24682 ;
  assign n33435 = ~n24684 ;
  assign n24685 = n24683 & n33435 ;
  assign n33436 = ~n24465 ;
  assign n24582 = n33436 & n24472 ;
  assign n24583 = n24464 | n24582 ;
  assign n33437 = ~n24435 ;
  assign n24584 = n33437 & n24442 ;
  assign n24585 = n24434 | n24584 ;
  assign n3879 = n1690 & n3876 ;
  assign n1608 = x[106] & n1551 ;
  assign n1630 = x[107] & n1616 ;
  assign n24586 = n1608 | n1630 ;
  assign n24587 = x[108] & n1547 ;
  assign n24588 = n24586 | n24587 ;
  assign n24589 = n3879 | n24588 ;
  assign n33438 = ~n24589 ;
  assign n24590 = x[53] & n33438 ;
  assign n24591 = n30125 & n24589 ;
  assign n24592 = n24590 | n24591 ;
  assign n33439 = ~n24418 ;
  assign n24593 = n24386 & n33439 ;
  assign n24594 = n24429 | n24593 ;
  assign n3411 = n1457 & n3409 ;
  assign n1339 = x[103] & n1319 ;
  assign n1401 = x[104] & n1384 ;
  assign n24595 = n1339 | n1401 ;
  assign n24596 = x[105] & n1315 ;
  assign n24597 = n24595 | n24596 ;
  assign n24598 = n3411 | n24597 ;
  assign n33440 = ~n24598 ;
  assign n24599 = x[56] & n33440 ;
  assign n24600 = n30379 & n24598 ;
  assign n24601 = n24599 | n24600 ;
  assign n33441 = ~n24403 ;
  assign n24404 = n24388 & n33441 ;
  assign n24602 = n24404 | n24415 ;
  assign n33442 = ~n24389 ;
  assign n24603 = n33442 & n24390 ;
  assign n33443 = ~n24393 ;
  assign n24604 = n33443 & n24400 ;
  assign n24605 = n24603 | n24604 ;
  assign n286 = x[95] & n27215 ;
  assign n828 = x[96] & n805 ;
  assign n24606 = n286 | n828 ;
  assign n33444 = ~n24606 ;
  assign n24607 = n24389 & n33444 ;
  assign n24608 = n33442 & n24606 ;
  assign n24609 = n24607 | n24608 ;
  assign n24610 = n24605 & n24609 ;
  assign n33445 = ~n24608 ;
  assign n24611 = n24605 & n33445 ;
  assign n24612 = n24607 | n24611 ;
  assign n24613 = n24608 | n24612 ;
  assign n33446 = ~n24610 ;
  assign n24614 = n33446 & n24613 ;
  assign n2320 = n1006 & n2313 ;
  assign n916 = x[97] & n900 ;
  assign n983 = x[98] & n949 ;
  assign n24615 = n916 | n983 ;
  assign n24616 = x[99] & n881 ;
  assign n24617 = n24615 | n24616 ;
  assign n24618 = n2320 | n24617 ;
  assign n33447 = ~n24618 ;
  assign n24619 = x[62] & n33447 ;
  assign n24620 = n30886 & n24618 ;
  assign n24621 = n24619 | n24620 ;
  assign n33448 = ~n24621 ;
  assign n24622 = n24614 & n33448 ;
  assign n33449 = ~n24614 ;
  assign n24623 = n33449 & n24621 ;
  assign n24624 = n24622 | n24623 ;
  assign n2875 = n1217 & n2867 ;
  assign n1109 = x[100] & n1079 ;
  assign n1196 = x[101] & n1144 ;
  assign n24625 = n1109 | n1196 ;
  assign n24626 = x[102] & n1075 ;
  assign n24627 = n24625 | n24626 ;
  assign n24628 = n2875 | n24627 ;
  assign n33450 = ~n24628 ;
  assign n24629 = x[59] & n33450 ;
  assign n24630 = n30638 & n24628 ;
  assign n24631 = n24629 | n24630 ;
  assign n24632 = n24624 & n24631 ;
  assign n24633 = n24624 | n24631 ;
  assign n33451 = ~n24632 ;
  assign n24634 = n33451 & n24633 ;
  assign n33452 = ~n24602 ;
  assign n24635 = n33452 & n24634 ;
  assign n33453 = ~n24634 ;
  assign n24636 = n24602 & n33453 ;
  assign n24637 = n24635 | n24636 ;
  assign n24638 = n24601 | n24637 ;
  assign n24640 = n24601 & n24637 ;
  assign n33454 = ~n24640 ;
  assign n24641 = n24638 & n33454 ;
  assign n24642 = n24594 | n24641 ;
  assign n24643 = n24594 & n24641 ;
  assign n33455 = ~n24643 ;
  assign n24644 = n24642 & n33455 ;
  assign n24645 = n24592 | n24644 ;
  assign n24646 = n24592 & n24644 ;
  assign n33456 = ~n24646 ;
  assign n24647 = n24645 & n33456 ;
  assign n24648 = n24585 | n24647 ;
  assign n24649 = n24585 & n24647 ;
  assign n33457 = ~n24649 ;
  assign n24650 = n24648 & n33457 ;
  assign n4254 = n2007 & n4246 ;
  assign n1883 = x[109] & n1866 ;
  assign n1985 = x[110] & n1931 ;
  assign n24651 = n1883 | n1985 ;
  assign n24652 = x[111] & n1862 ;
  assign n24653 = n24651 | n24652 ;
  assign n24654 = n4254 | n24653 ;
  assign n33458 = ~n24654 ;
  assign n24655 = x[50] & n33458 ;
  assign n24656 = n29865 & n24654 ;
  assign n24657 = n24655 | n24656 ;
  assign n24658 = n24650 | n24657 ;
  assign n24659 = n24650 & n24657 ;
  assign n33459 = ~n24659 ;
  assign n24660 = n24658 & n33459 ;
  assign n33460 = ~n24445 ;
  assign n24661 = n33460 & n24448 ;
  assign n33461 = ~n24451 ;
  assign n24662 = n33461 & n24458 ;
  assign n24663 = n24661 | n24662 ;
  assign n33462 = ~n24663 ;
  assign n24664 = n24660 & n33462 ;
  assign n33463 = ~n24660 ;
  assign n24665 = n33463 & n24663 ;
  assign n24666 = n24664 | n24665 ;
  assign n4280 = n2321 & n4276 ;
  assign n2212 = x[112] & n2179 ;
  assign n2262 = x[113] & n2244 ;
  assign n24667 = n2212 | n2262 ;
  assign n24668 = x[114] & n2175 ;
  assign n24669 = n24667 | n24668 ;
  assign n24670 = n4280 | n24669 ;
  assign n33464 = ~n24670 ;
  assign n24671 = x[47] & n33464 ;
  assign n24672 = n29621 & n24670 ;
  assign n24673 = n24671 | n24672 ;
  assign n24674 = n24666 | n24673 ;
  assign n24675 = n24666 & n24673 ;
  assign n33465 = ~n24675 ;
  assign n24676 = n24674 & n33465 ;
  assign n24677 = n24583 | n24676 ;
  assign n24678 = n24583 & n24676 ;
  assign n33466 = ~n24678 ;
  assign n24686 = n24677 & n33466 ;
  assign n33467 = ~n24686 ;
  assign n24687 = n24685 & n33467 ;
  assign n33468 = ~n24685 ;
  assign n24688 = n24677 & n33468 ;
  assign n24689 = n33466 & n24688 ;
  assign n24690 = n24687 | n24689 ;
  assign n33469 = ~n24581 ;
  assign n24691 = n33469 & n24690 ;
  assign n33470 = ~n24690 ;
  assign n24692 = n24581 & n33470 ;
  assign n24693 = n24691 | n24692 ;
  assign n24694 = n24579 | n24693 ;
  assign n24695 = n24579 & n24693 ;
  assign n33471 = ~n24695 ;
  assign n24696 = n24694 & n33471 ;
  assign n33472 = ~n24696 ;
  assign n24697 = n24572 & n33472 ;
  assign n33473 = ~n24572 ;
  assign n24698 = n33473 & n24696 ;
  assign n24699 = n24697 | n24698 ;
  assign n5418 = n3574 & n5417 ;
  assign n3445 = x[121] & n3443 ;
  assign n3551 = x[122] & n3508 ;
  assign n24700 = n3445 | n3551 ;
  assign n24701 = x[123] & n3439 ;
  assign n24702 = n24700 | n24701 ;
  assign n24703 = n5418 | n24702 ;
  assign n33474 = ~n24703 ;
  assign n24704 = x[38] & n33474 ;
  assign n24705 = n28996 & n24703 ;
  assign n24706 = n24704 | n24705 ;
  assign n24707 = n24699 | n24706 ;
  assign n24708 = n24699 & n24706 ;
  assign n33475 = ~n24708 ;
  assign n24709 = n24707 & n33475 ;
  assign n33476 = ~n24507 ;
  assign n24710 = n33476 & n24514 ;
  assign n24711 = n24505 | n24710 ;
  assign n33477 = ~n24711 ;
  assign n24712 = n24709 & n33477 ;
  assign n33478 = ~n24709 ;
  assign n24713 = n33478 & n24711 ;
  assign n24714 = n24712 | n24713 ;
  assign n5392 = n4041 & n5388 ;
  assign n3971 = x[124] & n3910 ;
  assign n3996 = x[125] & n3975 ;
  assign n24715 = n3971 | n3996 ;
  assign n24716 = x[126] & n3906 ;
  assign n24717 = n24715 | n24716 ;
  assign n24718 = n5392 | n24717 ;
  assign n33479 = ~n24718 ;
  assign n24719 = x[35] & n33479 ;
  assign n24720 = n28822 & n24718 ;
  assign n24721 = n24719 | n24720 ;
  assign n24722 = n24714 | n24721 ;
  assign n24723 = n24714 & n24721 ;
  assign n33480 = ~n24723 ;
  assign n24724 = n24722 & n33480 ;
  assign n33481 = ~n24570 ;
  assign n24725 = n33481 & n24724 ;
  assign n33482 = ~n24724 ;
  assign n24726 = n24570 & n33482 ;
  assign n24727 = n24725 | n24726 ;
  assign n24728 = n24562 & n24727 ;
  assign n24730 = n24562 | n24727 ;
  assign n33483 = ~n24728 ;
  assign n24731 = n33483 & n24730 ;
  assign n24732 = n24729 | n24731 ;
  assign n24733 = n24729 & n24730 ;
  assign n24734 = n33483 & n24733 ;
  assign n33484 = ~n24734 ;
  assign n224 = n24732 & n33484 ;
  assign n33485 = ~n24727 ;
  assign n24736 = n24562 & n33485 ;
  assign n33486 = ~n24736 ;
  assign n24737 = n24732 & n33486 ;
  assign n24738 = n24569 | n24726 ;
  assign n33487 = ~n24676 ;
  assign n24739 = n24583 & n33487 ;
  assign n24740 = n24687 | n24739 ;
  assign n33488 = ~n24666 ;
  assign n24741 = n33488 & n24673 ;
  assign n24742 = n24665 | n24741 ;
  assign n33489 = ~n24624 ;
  assign n24743 = n33489 & n24631 ;
  assign n24744 = n24623 | n24743 ;
  assign n287 = x[96] & n27215 ;
  assign n827 = x[97] & n805 ;
  assign n24745 = n287 | n827 ;
  assign n33490 = ~n24745 ;
  assign n24746 = x[32] & n33490 ;
  assign n24747 = n28658 & n24745 ;
  assign n24748 = n24746 | n24747 ;
  assign n24749 = n24606 | n24748 ;
  assign n24751 = n24606 & n24748 ;
  assign n33491 = ~n24751 ;
  assign n24752 = n24749 & n33491 ;
  assign n24753 = n24612 & n24752 ;
  assign n24754 = n24612 | n24752 ;
  assign n33492 = ~n24753 ;
  assign n24755 = n33492 & n24754 ;
  assign n2473 = n1006 & n2466 ;
  assign n903 = x[98] & n900 ;
  assign n954 = x[99] & n949 ;
  assign n24756 = n903 | n954 ;
  assign n24757 = x[100] & n881 ;
  assign n24758 = n24756 | n24757 ;
  assign n24759 = n2473 | n24758 ;
  assign n33493 = ~n24759 ;
  assign n24760 = x[62] & n33493 ;
  assign n24761 = n30886 & n24759 ;
  assign n24762 = n24760 | n24761 ;
  assign n33494 = ~n24762 ;
  assign n24763 = n24755 & n33494 ;
  assign n33495 = ~n24755 ;
  assign n24764 = n33495 & n24762 ;
  assign n24765 = n24763 | n24764 ;
  assign n2634 = n1217 & n2626 ;
  assign n1095 = x[101] & n1079 ;
  assign n1175 = x[102] & n1144 ;
  assign n24766 = n1095 | n1175 ;
  assign n24767 = x[103] & n1075 ;
  assign n24768 = n24766 | n24767 ;
  assign n24769 = n2634 | n24768 ;
  assign n33496 = ~n24769 ;
  assign n24770 = x[59] & n33496 ;
  assign n24771 = n30638 & n24769 ;
  assign n24772 = n24770 | n24771 ;
  assign n33497 = ~n24772 ;
  assign n24773 = n24765 & n33497 ;
  assign n33498 = ~n24765 ;
  assign n24774 = n33498 & n24772 ;
  assign n24775 = n24773 | n24774 ;
  assign n24776 = n24744 | n24775 ;
  assign n24777 = n24744 & n24775 ;
  assign n33499 = ~n24777 ;
  assign n24778 = n24776 & n33499 ;
  assign n3231 = n1457 & n3223 ;
  assign n1338 = x[104] & n1319 ;
  assign n1399 = x[105] & n1384 ;
  assign n24779 = n1338 | n1399 ;
  assign n24780 = x[106] & n1315 ;
  assign n24781 = n24779 | n24780 ;
  assign n24782 = n3231 | n24781 ;
  assign n33500 = ~n24782 ;
  assign n24783 = x[56] & n33500 ;
  assign n24784 = n30379 & n24782 ;
  assign n24785 = n24783 | n24784 ;
  assign n24786 = n24778 | n24785 ;
  assign n24787 = n24778 & n24785 ;
  assign n33501 = ~n24787 ;
  assign n24788 = n24786 & n33501 ;
  assign n33502 = ~n24637 ;
  assign n24639 = n24601 & n33502 ;
  assign n24789 = n24636 | n24639 ;
  assign n24790 = n24788 | n24789 ;
  assign n24791 = n24788 & n24789 ;
  assign n33503 = ~n24791 ;
  assign n24792 = n24790 & n33503 ;
  assign n3648 = n1690 & n3639 ;
  assign n1560 = x[107] & n1551 ;
  assign n1626 = x[108] & n1616 ;
  assign n24793 = n1560 | n1626 ;
  assign n24794 = x[109] & n1547 ;
  assign n24795 = n24793 | n24794 ;
  assign n24796 = n3648 | n24795 ;
  assign n33504 = ~n24796 ;
  assign n24797 = x[53] & n33504 ;
  assign n24798 = n30125 & n24796 ;
  assign n24799 = n24797 | n24798 ;
  assign n24800 = n24792 | n24799 ;
  assign n24801 = n24792 & n24799 ;
  assign n33505 = ~n24801 ;
  assign n24802 = n24800 & n33505 ;
  assign n33506 = ~n24641 ;
  assign n24803 = n24594 & n33506 ;
  assign n33507 = ~n24644 ;
  assign n24804 = n24592 & n33507 ;
  assign n24805 = n24803 | n24804 ;
  assign n24806 = n24802 | n24805 ;
  assign n24807 = n24802 & n24805 ;
  assign n33508 = ~n24807 ;
  assign n24808 = n24806 & n33508 ;
  assign n4450 = n2007 & n4442 ;
  assign n1890 = x[110] & n1866 ;
  assign n1939 = x[111] & n1931 ;
  assign n24809 = n1890 | n1939 ;
  assign n24810 = x[112] & n1862 ;
  assign n24811 = n24809 | n24810 ;
  assign n24812 = n4450 | n24811 ;
  assign n33509 = ~n24812 ;
  assign n24813 = x[50] & n33509 ;
  assign n24814 = n29865 & n24812 ;
  assign n24815 = n24813 | n24814 ;
  assign n24816 = n24808 | n24815 ;
  assign n24817 = n24808 & n24815 ;
  assign n33510 = ~n24817 ;
  assign n24818 = n24816 & n33510 ;
  assign n33511 = ~n24647 ;
  assign n24819 = n24585 & n33511 ;
  assign n33512 = ~n24650 ;
  assign n24820 = n33512 & n24657 ;
  assign n24821 = n24819 | n24820 ;
  assign n24822 = n24818 | n24821 ;
  assign n24823 = n24818 & n24821 ;
  assign n33513 = ~n24823 ;
  assign n24824 = n24822 & n33513 ;
  assign n4478 = n2321 & n4474 ;
  assign n2192 = x[113] & n2179 ;
  assign n2252 = x[114] & n2244 ;
  assign n24825 = n2192 | n2252 ;
  assign n24826 = x[115] & n2175 ;
  assign n24827 = n24825 | n24826 ;
  assign n24828 = n4478 | n24827 ;
  assign n33514 = ~n24828 ;
  assign n24829 = x[47] & n33514 ;
  assign n24830 = n29621 & n24828 ;
  assign n24831 = n24829 | n24830 ;
  assign n33515 = ~n24824 ;
  assign n24832 = n33515 & n24831 ;
  assign n33516 = ~n24831 ;
  assign n24833 = n24824 & n33516 ;
  assign n24834 = n24832 | n24833 ;
  assign n24835 = n24742 & n24834 ;
  assign n33517 = ~n24833 ;
  assign n24836 = n24742 & n33517 ;
  assign n24837 = n24832 | n24836 ;
  assign n24838 = n24833 | n24837 ;
  assign n33518 = ~n24835 ;
  assign n24839 = n33518 & n24838 ;
  assign n2646 = n784 & n2635 ;
  assign n2544 = x[116] & n2492 ;
  assign n2574 = x[117] & n2557 ;
  assign n24840 = n2544 | n2574 ;
  assign n24841 = x[118] & n2488 ;
  assign n24842 = n24840 | n24841 ;
  assign n24843 = n2646 | n24842 ;
  assign n33519 = ~n24843 ;
  assign n24844 = x[44] & n33519 ;
  assign n24845 = n29400 & n24843 ;
  assign n24846 = n24844 | n24845 ;
  assign n33520 = ~n24846 ;
  assign n24847 = n24839 & n33520 ;
  assign n33521 = ~n24839 ;
  assign n24848 = n33521 & n24846 ;
  assign n24849 = n24847 | n24848 ;
  assign n24850 = n24740 | n24849 ;
  assign n24851 = n24740 & n24849 ;
  assign n33522 = ~n24851 ;
  assign n24852 = n24850 & n33522 ;
  assign n4993 = n3162 & n4985 ;
  assign n3080 = x[119] & n3031 ;
  assign n3099 = x[120] & n3096 ;
  assign n24853 = n3080 | n3099 ;
  assign n24854 = x[121] & n3027 ;
  assign n24855 = n24853 | n24854 ;
  assign n24856 = n4993 | n24855 ;
  assign n33523 = ~n24856 ;
  assign n24857 = x[41] & n33523 ;
  assign n24858 = n29184 & n24856 ;
  assign n24859 = n24857 | n24858 ;
  assign n24860 = n24852 | n24859 ;
  assign n24861 = n24852 & n24859 ;
  assign n33524 = ~n24861 ;
  assign n24862 = n24860 & n33524 ;
  assign n33525 = ~n24693 ;
  assign n24863 = n24579 & n33525 ;
  assign n24864 = n24692 | n24863 ;
  assign n24865 = n24862 | n24864 ;
  assign n24866 = n24862 & n24864 ;
  assign n33526 = ~n24866 ;
  assign n24867 = n24865 & n33526 ;
  assign n5841 = n3574 & n5838 ;
  assign n3444 = x[122] & n3443 ;
  assign n3550 = x[123] & n3508 ;
  assign n24868 = n3444 | n3550 ;
  assign n24869 = x[124] & n3439 ;
  assign n24870 = n24868 | n24869 ;
  assign n24871 = n5841 | n24870 ;
  assign n33527 = ~n24871 ;
  assign n24872 = x[38] & n33527 ;
  assign n24873 = n28996 & n24871 ;
  assign n24874 = n24872 | n24873 ;
  assign n24875 = n24867 | n24874 ;
  assign n24876 = n24867 & n24874 ;
  assign n33528 = ~n24876 ;
  assign n24877 = n24875 & n33528 ;
  assign n33529 = ~n24699 ;
  assign n24878 = n33529 & n24706 ;
  assign n24879 = n24697 | n24878 ;
  assign n33530 = ~n24879 ;
  assign n24880 = n24877 & n33530 ;
  assign n33531 = ~n24877 ;
  assign n24881 = n33531 & n24879 ;
  assign n24882 = n24880 | n24881 ;
  assign n33532 = ~n24714 ;
  assign n24883 = n33532 & n24721 ;
  assign n24884 = n24713 | n24883 ;
  assign n5630 = n4041 & n5629 ;
  assign n3972 = x[125] & n3910 ;
  assign n4028 = x[126] & n3975 ;
  assign n24885 = n3972 | n4028 ;
  assign n24886 = x[127] & n3906 ;
  assign n24887 = n24885 | n24886 ;
  assign n24888 = n5630 | n24887 ;
  assign n33533 = ~n24888 ;
  assign n24889 = x[35] & n33533 ;
  assign n24890 = n28822 & n24888 ;
  assign n24891 = n24889 | n24890 ;
  assign n33534 = ~n24891 ;
  assign n24892 = n24884 & n33534 ;
  assign n33535 = ~n24884 ;
  assign n24893 = n33535 & n24891 ;
  assign n24894 = n24892 | n24893 ;
  assign n24895 = n24882 | n24894 ;
  assign n24896 = n24882 & n24894 ;
  assign n33536 = ~n24896 ;
  assign n24897 = n24895 & n33536 ;
  assign n33537 = ~n24897 ;
  assign n24898 = n24738 & n33537 ;
  assign n33538 = ~n24738 ;
  assign n24899 = n33538 & n24897 ;
  assign n24900 = n24898 | n24899 ;
  assign n24901 = n24737 | n24900 ;
  assign n24902 = n24737 & n24900 ;
  assign n33539 = ~n24902 ;
  assign n225 = n24901 & n33539 ;
  assign n33540 = ~n24867 ;
  assign n25041 = n33540 & n24874 ;
  assign n25042 = n24881 | n25041 ;
  assign n6187 = n4041 & n6186 ;
  assign n3973 = x[126] & n3910 ;
  assign n25043 = x[127] & n3975 ;
  assign n25044 = n3973 | n25043 ;
  assign n25045 = n6187 | n25044 ;
  assign n33541 = ~n25045 ;
  assign n25046 = x[35] & n33541 ;
  assign n25047 = n28822 & n25045 ;
  assign n25048 = n25046 | n25047 ;
  assign n25049 = n25042 | n25048 ;
  assign n25050 = n25042 & n25048 ;
  assign n33542 = ~n25050 ;
  assign n25051 = n25049 & n33542 ;
  assign n33543 = ~n24849 ;
  assign n24904 = n24740 & n33543 ;
  assign n24905 = n24848 | n24904 ;
  assign n33544 = ~n24775 ;
  assign n24906 = n24744 & n33544 ;
  assign n24907 = n24774 | n24906 ;
  assign n3003 = n1217 & n3001 ;
  assign n1094 = x[102] & n1079 ;
  assign n1158 = x[103] & n1144 ;
  assign n24927 = n1094 | n1158 ;
  assign n24928 = x[104] & n1075 ;
  assign n24929 = n24927 | n24928 ;
  assign n24930 = n3003 | n24929 ;
  assign n24931 = x[59] | n24930 ;
  assign n24932 = x[59] & n24930 ;
  assign n33545 = ~n24932 ;
  assign n24933 = n24931 & n33545 ;
  assign n33546 = ~n24752 ;
  assign n24908 = n24612 & n33546 ;
  assign n24909 = n24764 | n24908 ;
  assign n288 = x[97] & n27215 ;
  assign n825 = x[98] & n805 ;
  assign n24910 = n288 | n825 ;
  assign n33547 = ~n24748 ;
  assign n24750 = n24606 & n33547 ;
  assign n24911 = n24747 | n24750 ;
  assign n24912 = n24910 | n24911 ;
  assign n24913 = n24910 & n24911 ;
  assign n33548 = ~n24913 ;
  assign n24914 = n24912 & n33548 ;
  assign n2981 = n1006 & n2977 ;
  assign n901 = x[99] & n900 ;
  assign n963 = x[100] & n949 ;
  assign n24915 = n901 | n963 ;
  assign n24916 = x[101] & n881 ;
  assign n24917 = n24915 | n24916 ;
  assign n24918 = n2981 | n24917 ;
  assign n33549 = ~n24918 ;
  assign n24919 = x[62] & n33549 ;
  assign n24920 = n30886 & n24918 ;
  assign n24921 = n24919 | n24920 ;
  assign n24922 = n24914 | n24921 ;
  assign n24923 = n24914 & n24921 ;
  assign n33550 = ~n24923 ;
  assign n24924 = n24922 & n33550 ;
  assign n24926 = n24909 & n24924 ;
  assign n24934 = n24909 | n24924 ;
  assign n33551 = ~n24926 ;
  assign n24935 = n33551 & n24934 ;
  assign n33552 = ~n24935 ;
  assign n24936 = n24933 & n33552 ;
  assign n33553 = ~n24933 ;
  assign n24937 = n33553 & n24934 ;
  assign n24938 = n33551 & n24937 ;
  assign n24939 = n24936 | n24938 ;
  assign n33554 = ~n24907 ;
  assign n24940 = n33554 & n24939 ;
  assign n33555 = ~n24939 ;
  assign n24941 = n24907 & n33555 ;
  assign n24942 = n24940 | n24941 ;
  assign n3201 = n1457 & n3199 ;
  assign n1336 = x[105] & n1319 ;
  assign n1402 = x[106] & n1384 ;
  assign n24943 = n1336 | n1402 ;
  assign n24944 = x[107] & n1315 ;
  assign n24945 = n24943 | n24944 ;
  assign n24946 = n3201 | n24945 ;
  assign n33556 = ~n24946 ;
  assign n24947 = x[56] & n33556 ;
  assign n24948 = n30379 & n24946 ;
  assign n24949 = n24947 | n24948 ;
  assign n24950 = n24942 | n24949 ;
  assign n24951 = n24942 & n24949 ;
  assign n33557 = ~n24951 ;
  assign n24952 = n24950 & n33557 ;
  assign n33558 = ~n24778 ;
  assign n24953 = n33558 & n24785 ;
  assign n33559 = ~n24788 ;
  assign n24954 = n33559 & n24789 ;
  assign n24955 = n24953 | n24954 ;
  assign n24956 = n24952 | n24955 ;
  assign n24957 = n24952 & n24955 ;
  assign n33560 = ~n24957 ;
  assign n24958 = n24956 & n33560 ;
  assign n3621 = n1690 & n3615 ;
  assign n1605 = x[108] & n1551 ;
  assign n1637 = x[109] & n1616 ;
  assign n24959 = n1605 | n1637 ;
  assign n24960 = x[110] & n1547 ;
  assign n24961 = n24959 | n24960 ;
  assign n24962 = n3621 | n24961 ;
  assign n33561 = ~n24962 ;
  assign n24963 = x[53] & n33561 ;
  assign n24964 = n30125 & n24962 ;
  assign n24965 = n24963 | n24964 ;
  assign n24966 = n24958 | n24965 ;
  assign n24967 = n24958 & n24965 ;
  assign n33562 = ~n24967 ;
  assign n24968 = n24966 & n33562 ;
  assign n33563 = ~n24792 ;
  assign n24969 = n33563 & n24799 ;
  assign n33564 = ~n24802 ;
  assign n24970 = n33564 & n24805 ;
  assign n24971 = n24969 | n24970 ;
  assign n33565 = ~n24971 ;
  assign n24972 = n24968 & n33565 ;
  assign n33566 = ~n24968 ;
  assign n24973 = n33566 & n24971 ;
  assign n24974 = n24972 | n24973 ;
  assign n4096 = n2007 & n4087 ;
  assign n1881 = x[111] & n1866 ;
  assign n1938 = x[112] & n1931 ;
  assign n24975 = n1881 | n1938 ;
  assign n24976 = x[113] & n1862 ;
  assign n24977 = n24975 | n24976 ;
  assign n24978 = n4096 | n24977 ;
  assign n33567 = ~n24978 ;
  assign n24979 = x[50] & n33567 ;
  assign n24980 = n29865 & n24978 ;
  assign n24981 = n24979 | n24980 ;
  assign n24982 = n24974 | n24981 ;
  assign n24983 = n24974 & n24981 ;
  assign n33568 = ~n24983 ;
  assign n24984 = n24982 & n33568 ;
  assign n33569 = ~n24808 ;
  assign n24985 = n33569 & n24815 ;
  assign n33570 = ~n24818 ;
  assign n24986 = n33570 & n24821 ;
  assign n24987 = n24985 | n24986 ;
  assign n33571 = ~n24987 ;
  assign n24988 = n24984 & n33571 ;
  assign n33572 = ~n24984 ;
  assign n24989 = n33572 & n24987 ;
  assign n24990 = n24988 | n24989 ;
  assign n4705 = n2321 & n4702 ;
  assign n2233 = x[114] & n2179 ;
  assign n2267 = x[115] & n2244 ;
  assign n24991 = n2233 | n2267 ;
  assign n24992 = x[116] & n2175 ;
  assign n24993 = n24991 | n24992 ;
  assign n24994 = n4705 | n24993 ;
  assign n33573 = ~n24994 ;
  assign n24995 = x[47] & n33573 ;
  assign n24996 = n29621 & n24994 ;
  assign n24997 = n24995 | n24996 ;
  assign n24998 = n24990 | n24997 ;
  assign n24999 = n24990 & n24997 ;
  assign n33574 = ~n24999 ;
  assign n25000 = n24998 & n33574 ;
  assign n25001 = n24837 & n25000 ;
  assign n25002 = n24837 | n25000 ;
  assign n33575 = ~n25001 ;
  assign n25003 = n33575 & n25002 ;
  assign n5056 = n2635 & n5047 ;
  assign n2502 = x[117] & n2492 ;
  assign n2581 = x[118] & n2557 ;
  assign n25004 = n2502 | n2581 ;
  assign n25005 = x[119] & n2488 ;
  assign n25006 = n25004 | n25005 ;
  assign n25007 = n5056 | n25006 ;
  assign n33576 = ~n25007 ;
  assign n25008 = x[44] & n33576 ;
  assign n25009 = n29400 & n25007 ;
  assign n25010 = n25008 | n25009 ;
  assign n33577 = ~n25010 ;
  assign n25011 = n25003 & n33577 ;
  assign n33578 = ~n25003 ;
  assign n25012 = n33578 & n25010 ;
  assign n25013 = n25011 | n25012 ;
  assign n33579 = ~n25013 ;
  assign n25014 = n24905 & n33579 ;
  assign n33580 = ~n24905 ;
  assign n25015 = n33580 & n25013 ;
  assign n25016 = n25014 | n25015 ;
  assign n5032 = n3162 & n5022 ;
  assign n3034 = x[120] & n3031 ;
  assign n3098 = x[121] & n3096 ;
  assign n25017 = n3034 | n3098 ;
  assign n25018 = x[122] & n3027 ;
  assign n25019 = n25017 | n25018 ;
  assign n25020 = n5032 | n25019 ;
  assign n33581 = ~n25020 ;
  assign n25021 = x[41] & n33581 ;
  assign n25022 = n29184 & n25020 ;
  assign n25023 = n25021 | n25022 ;
  assign n25024 = n25016 | n25023 ;
  assign n25025 = n25016 & n25023 ;
  assign n33582 = ~n25025 ;
  assign n25026 = n25024 & n33582 ;
  assign n33583 = ~n24852 ;
  assign n25027 = n33583 & n24859 ;
  assign n33584 = ~n24862 ;
  assign n25028 = n33584 & n24864 ;
  assign n25029 = n25027 | n25028 ;
  assign n33585 = ~n25029 ;
  assign n25030 = n25026 & n33585 ;
  assign n33586 = ~n25026 ;
  assign n25031 = n33586 & n25029 ;
  assign n25032 = n25030 | n25031 ;
  assign n3611 = n642 & n3574 ;
  assign n3506 = x[123] & n3443 ;
  assign n3569 = x[124] & n3508 ;
  assign n25033 = n3506 | n3569 ;
  assign n25034 = x[125] & n3439 ;
  assign n25035 = n25033 | n25034 ;
  assign n25036 = n3611 | n25035 ;
  assign n33587 = ~n25036 ;
  assign n25037 = x[38] & n33587 ;
  assign n25038 = n28996 & n25036 ;
  assign n25039 = n25037 | n25038 ;
  assign n33588 = ~n25032 ;
  assign n25040 = n33588 & n25039 ;
  assign n33589 = ~n25039 ;
  assign n25052 = n25032 & n33589 ;
  assign n33590 = ~n25052 ;
  assign n25053 = n25051 & n33590 ;
  assign n33591 = ~n25040 ;
  assign n25054 = n33591 & n25053 ;
  assign n33592 = ~n25054 ;
  assign n25055 = n25051 & n33592 ;
  assign n25056 = n25052 | n25054 ;
  assign n25057 = n25040 | n25056 ;
  assign n33593 = ~n25055 ;
  assign n25058 = n33593 & n25057 ;
  assign n25059 = n24884 & n24891 ;
  assign n33594 = ~n24882 ;
  assign n25060 = n33594 & n24894 ;
  assign n25061 = n25059 | n25060 ;
  assign n33595 = ~n25061 ;
  assign n25062 = n25058 & n33595 ;
  assign n33596 = ~n25058 ;
  assign n25063 = n33596 & n25061 ;
  assign n25064 = n25062 | n25063 ;
  assign n33597 = ~n24898 ;
  assign n25065 = n33597 & n24901 ;
  assign n25066 = n25064 & n25065 ;
  assign n25067 = n25064 | n25065 ;
  assign n33598 = ~n25066 ;
  assign n226 = n33598 & n25067 ;
  assign n33599 = ~n25063 ;
  assign n25069 = n33599 & n25067 ;
  assign n25070 = n25050 | n25054 ;
  assign n25071 = n25031 | n25040 ;
  assign n3974 = x[127] & n3910 ;
  assign n5366 = n4041 & n5360 ;
  assign n25072 = n3974 | n5366 ;
  assign n33600 = ~n25072 ;
  assign n25073 = x[35] & n33600 ;
  assign n25074 = n28822 & n25072 ;
  assign n25075 = n25073 | n25074 ;
  assign n25076 = n25071 | n25075 ;
  assign n25077 = n25071 & n25075 ;
  assign n33601 = ~n25077 ;
  assign n25078 = n25076 & n33601 ;
  assign n33602 = ~n25000 ;
  assign n25079 = n24837 & n33602 ;
  assign n25080 = n25012 | n25079 ;
  assign n4681 = n2635 & n4678 ;
  assign n2511 = x[118] & n2492 ;
  assign n2577 = x[119] & n2557 ;
  assign n25081 = n2511 | n2577 ;
  assign n25082 = x[120] & n2488 ;
  assign n25083 = n25081 | n25082 ;
  assign n25084 = n4681 | n25083 ;
  assign n33603 = ~n25084 ;
  assign n25085 = x[44] & n33603 ;
  assign n25086 = n29400 & n25084 ;
  assign n25087 = n25085 | n25086 ;
  assign n33604 = ~n24990 ;
  assign n25088 = n33604 & n24997 ;
  assign n25089 = n24989 | n25088 ;
  assign n2322 = n797 & n2321 ;
  assign n2182 = x[115] & n2179 ;
  assign n2250 = x[116] & n2244 ;
  assign n25173 = n2182 | n2250 ;
  assign n25174 = x[117] & n2175 ;
  assign n25175 = n25173 | n25174 ;
  assign n25176 = n2322 | n25175 ;
  assign n25177 = x[47] | n25176 ;
  assign n25178 = x[47] & n25176 ;
  assign n33605 = ~n25178 ;
  assign n25179 = n25177 & n33605 ;
  assign n33606 = ~n24974 ;
  assign n25090 = n33606 & n24981 ;
  assign n25091 = n24973 | n25090 ;
  assign n33607 = ~n24942 ;
  assign n25092 = n33607 & n24949 ;
  assign n25093 = n24941 | n25092 ;
  assign n3883 = n1457 & n3876 ;
  assign n1335 = x[106] & n1319 ;
  assign n1397 = x[107] & n1384 ;
  assign n25094 = n1335 | n1397 ;
  assign n25095 = x[108] & n1315 ;
  assign n25096 = n25094 | n25095 ;
  assign n25097 = n3883 | n25096 ;
  assign n33608 = ~n25097 ;
  assign n25098 = x[56] & n33608 ;
  assign n25099 = n30379 & n25097 ;
  assign n25100 = n25098 | n25099 ;
  assign n33609 = ~n24924 ;
  assign n24925 = n24909 & n33609 ;
  assign n25101 = n24925 | n24936 ;
  assign n33610 = ~n24910 ;
  assign n25105 = n33610 & n24911 ;
  assign n33611 = ~n24914 ;
  assign n25106 = n33611 & n24921 ;
  assign n25108 = n25105 | n25106 ;
  assign n289 = x[98] & n27215 ;
  assign n823 = x[99] & n805 ;
  assign n25102 = n289 | n823 ;
  assign n25104 = n33610 & n25102 ;
  assign n33612 = ~n25102 ;
  assign n25107 = n24910 & n33612 ;
  assign n25109 = n25104 | n25107 ;
  assign n25110 = n25108 & n25109 ;
  assign n33613 = ~n25104 ;
  assign n25111 = n33613 & n25108 ;
  assign n25112 = n25107 | n25111 ;
  assign n25113 = n25104 | n25112 ;
  assign n33614 = ~n25110 ;
  assign n25114 = n33614 & n25113 ;
  assign n2869 = n1006 & n2867 ;
  assign n913 = x[100] & n900 ;
  assign n950 = x[101] & n949 ;
  assign n25115 = n913 | n950 ;
  assign n25116 = x[102] & n881 ;
  assign n25117 = n25115 | n25116 ;
  assign n25118 = n2869 | n25117 ;
  assign n33615 = ~n25118 ;
  assign n25119 = x[62] & n33615 ;
  assign n25120 = n30886 & n25118 ;
  assign n25121 = n25119 | n25120 ;
  assign n25122 = n25114 | n25121 ;
  assign n25123 = n25114 & n25121 ;
  assign n33616 = ~n25123 ;
  assign n25124 = n25122 & n33616 ;
  assign n3412 = n1217 & n3409 ;
  assign n1086 = x[103] & n1079 ;
  assign n1168 = x[104] & n1144 ;
  assign n25125 = n1086 | n1168 ;
  assign n25126 = x[105] & n1075 ;
  assign n25127 = n25125 | n25126 ;
  assign n25128 = n3412 | n25127 ;
  assign n33617 = ~n25128 ;
  assign n25129 = x[59] & n33617 ;
  assign n25130 = n30638 & n25128 ;
  assign n25131 = n25129 | n25130 ;
  assign n25133 = n25124 | n25131 ;
  assign n25134 = n25124 & n25131 ;
  assign n33618 = ~n25134 ;
  assign n25135 = n25133 & n33618 ;
  assign n33619 = ~n25101 ;
  assign n25136 = n33619 & n25135 ;
  assign n33620 = ~n25135 ;
  assign n25137 = n25101 & n33620 ;
  assign n25138 = n25136 | n25137 ;
  assign n25139 = n25100 | n25138 ;
  assign n25140 = n25100 & n25138 ;
  assign n33621 = ~n25140 ;
  assign n25141 = n25139 & n33621 ;
  assign n25142 = n25093 | n25141 ;
  assign n25143 = n25093 & n25141 ;
  assign n33622 = ~n25143 ;
  assign n25144 = n25142 & n33622 ;
  assign n4255 = n1690 & n4246 ;
  assign n1578 = x[109] & n1551 ;
  assign n1629 = x[110] & n1616 ;
  assign n25145 = n1578 | n1629 ;
  assign n25146 = x[111] & n1547 ;
  assign n25147 = n25145 | n25146 ;
  assign n25148 = n4255 | n25147 ;
  assign n33623 = ~n25148 ;
  assign n25149 = x[53] & n33623 ;
  assign n25150 = n30125 & n25148 ;
  assign n25151 = n25149 | n25150 ;
  assign n25152 = n25144 | n25151 ;
  assign n25153 = n25144 & n25151 ;
  assign n33624 = ~n25153 ;
  assign n25154 = n25152 & n33624 ;
  assign n33625 = ~n24952 ;
  assign n25155 = n33625 & n24955 ;
  assign n33626 = ~n24958 ;
  assign n25156 = n33626 & n24965 ;
  assign n25157 = n25155 | n25156 ;
  assign n33627 = ~n25157 ;
  assign n25158 = n25154 & n33627 ;
  assign n33628 = ~n25154 ;
  assign n25159 = n33628 & n25157 ;
  assign n25160 = n25158 | n25159 ;
  assign n4284 = n2007 & n4276 ;
  assign n1878 = x[112] & n1866 ;
  assign n1974 = x[113] & n1931 ;
  assign n25161 = n1878 | n1974 ;
  assign n25162 = x[114] & n1862 ;
  assign n25163 = n25161 | n25162 ;
  assign n25164 = n4284 | n25163 ;
  assign n33629 = ~n25164 ;
  assign n25165 = x[50] & n33629 ;
  assign n25166 = n29865 & n25164 ;
  assign n25167 = n25165 | n25166 ;
  assign n25168 = n25160 | n25167 ;
  assign n25169 = n25160 & n25167 ;
  assign n33630 = ~n25169 ;
  assign n25170 = n25168 & n33630 ;
  assign n25171 = n25091 | n25170 ;
  assign n25172 = n25091 & n25170 ;
  assign n33631 = ~n25172 ;
  assign n25180 = n25171 & n33631 ;
  assign n33632 = ~n25180 ;
  assign n25181 = n25179 & n33632 ;
  assign n33633 = ~n25179 ;
  assign n25182 = n25171 & n33633 ;
  assign n25183 = n33631 & n25182 ;
  assign n25184 = n25181 | n25183 ;
  assign n33634 = ~n25089 ;
  assign n25185 = n33634 & n25184 ;
  assign n33635 = ~n25184 ;
  assign n25186 = n25089 & n33635 ;
  assign n25187 = n25185 | n25186 ;
  assign n25188 = n25087 | n25187 ;
  assign n25189 = n25087 & n25187 ;
  assign n33636 = ~n25189 ;
  assign n25190 = n25188 & n33636 ;
  assign n33637 = ~n25190 ;
  assign n25191 = n25080 & n33637 ;
  assign n33638 = ~n25080 ;
  assign n25192 = n33638 & n25190 ;
  assign n25193 = n25191 | n25192 ;
  assign n5427 = n3162 & n5417 ;
  assign n3058 = x[121] & n3031 ;
  assign n3097 = x[122] & n3096 ;
  assign n25194 = n3058 | n3097 ;
  assign n25195 = x[123] & n3027 ;
  assign n25196 = n25194 | n25195 ;
  assign n25197 = n5427 | n25196 ;
  assign n33639 = ~n25197 ;
  assign n25198 = x[41] & n33639 ;
  assign n25199 = n29184 & n25197 ;
  assign n25200 = n25198 | n25199 ;
  assign n25201 = n25193 | n25200 ;
  assign n25202 = n25193 & n25200 ;
  assign n33640 = ~n25202 ;
  assign n25203 = n25201 & n33640 ;
  assign n33641 = ~n25016 ;
  assign n25204 = n33641 & n25023 ;
  assign n25205 = n25014 | n25204 ;
  assign n33642 = ~n25205 ;
  assign n25206 = n25203 & n33642 ;
  assign n33643 = ~n25203 ;
  assign n25207 = n33643 & n25205 ;
  assign n25208 = n25206 | n25207 ;
  assign n5396 = n3574 & n5388 ;
  assign n3448 = x[124] & n3443 ;
  assign n3570 = x[125] & n3508 ;
  assign n25209 = n3448 | n3570 ;
  assign n25210 = x[126] & n3439 ;
  assign n25211 = n25209 | n25210 ;
  assign n25212 = n5396 | n25211 ;
  assign n33644 = ~n25212 ;
  assign n25213 = x[38] & n33644 ;
  assign n25214 = n28996 & n25212 ;
  assign n25215 = n25213 | n25214 ;
  assign n25216 = n25208 | n25215 ;
  assign n25217 = n25208 & n25215 ;
  assign n33645 = ~n25217 ;
  assign n25218 = n25216 & n33645 ;
  assign n25220 = n25078 & n25218 ;
  assign n25221 = n25078 | n25218 ;
  assign n33646 = ~n25220 ;
  assign n25222 = n33646 & n25221 ;
  assign n33647 = ~n25070 ;
  assign n25223 = n33647 & n25222 ;
  assign n33648 = ~n25222 ;
  assign n25224 = n25070 & n33648 ;
  assign n25225 = n25223 | n25224 ;
  assign n25226 = n25069 | n25225 ;
  assign n25227 = n25069 & n25225 ;
  assign n33649 = ~n25227 ;
  assign n227 = n25226 & n33649 ;
  assign n33650 = ~n25224 ;
  assign n25229 = n33650 & n25226 ;
  assign n33651 = ~n25170 ;
  assign n25230 = n25091 & n33651 ;
  assign n25231 = n25181 | n25230 ;
  assign n2332 = n784 & n2321 ;
  assign n2186 = x[116] & n2179 ;
  assign n2249 = x[117] & n2244 ;
  assign n25232 = n2186 | n2249 ;
  assign n25233 = x[118] & n2175 ;
  assign n25234 = n25232 | n25233 ;
  assign n25235 = n2332 | n25234 ;
  assign n25236 = x[47] | n25235 ;
  assign n25237 = x[47] & n25235 ;
  assign n33652 = ~n25237 ;
  assign n25238 = n25236 & n33652 ;
  assign n33653 = ~n25160 ;
  assign n25239 = n33653 & n25167 ;
  assign n25240 = n25159 | n25239 ;
  assign n290 = x[99] & n27215 ;
  assign n822 = x[100] & n805 ;
  assign n25241 = n290 | n822 ;
  assign n25103 = x[35] | n25102 ;
  assign n25242 = x[35] & n25102 ;
  assign n33654 = ~n25242 ;
  assign n25243 = n25103 & n33654 ;
  assign n33655 = ~n25241 ;
  assign n25244 = n33655 & n25243 ;
  assign n33656 = ~n25243 ;
  assign n25245 = n25241 & n33656 ;
  assign n25246 = n25244 | n25245 ;
  assign n33657 = ~n25246 ;
  assign n25247 = n25112 & n33657 ;
  assign n33658 = ~n25112 ;
  assign n25248 = n33658 & n25246 ;
  assign n25249 = n25247 | n25248 ;
  assign n2630 = n1006 & n2626 ;
  assign n902 = x[101] & n900 ;
  assign n989 = x[102] & n949 ;
  assign n25250 = n902 | n989 ;
  assign n25251 = x[103] & n881 ;
  assign n25252 = n25250 | n25251 ;
  assign n25253 = n2630 | n25252 ;
  assign n33659 = ~n25253 ;
  assign n25254 = x[62] & n33659 ;
  assign n25255 = n30886 & n25253 ;
  assign n25256 = n25254 | n25255 ;
  assign n25257 = n25249 | n25256 ;
  assign n25258 = n25249 & n25256 ;
  assign n33660 = ~n25258 ;
  assign n25259 = n25257 & n33660 ;
  assign n3233 = n1217 & n3223 ;
  assign n1123 = x[104] & n1079 ;
  assign n1157 = x[105] & n1144 ;
  assign n25260 = n1123 | n1157 ;
  assign n25261 = x[106] & n1075 ;
  assign n25262 = n25260 | n25261 ;
  assign n25263 = n3233 | n25262 ;
  assign n33661 = ~n25263 ;
  assign n25264 = x[59] & n33661 ;
  assign n25265 = n30638 & n25263 ;
  assign n25266 = n25264 | n25265 ;
  assign n25267 = n25259 | n25266 ;
  assign n25268 = n25259 & n25266 ;
  assign n33662 = ~n25268 ;
  assign n25269 = n25267 & n33662 ;
  assign n33663 = ~n25124 ;
  assign n25132 = n33663 & n25131 ;
  assign n33664 = ~n25114 ;
  assign n25270 = n33664 & n25121 ;
  assign n25271 = n25132 | n25270 ;
  assign n33665 = ~n25271 ;
  assign n25272 = n25269 & n33665 ;
  assign n33666 = ~n25269 ;
  assign n25273 = n33666 & n25271 ;
  assign n25274 = n25272 | n25273 ;
  assign n3642 = n1457 & n3639 ;
  assign n1333 = x[107] & n1319 ;
  assign n1426 = x[108] & n1384 ;
  assign n25275 = n1333 | n1426 ;
  assign n25276 = x[109] & n1315 ;
  assign n25277 = n25275 | n25276 ;
  assign n25278 = n3642 | n25277 ;
  assign n33667 = ~n25278 ;
  assign n25279 = x[56] & n33667 ;
  assign n25280 = n30379 & n25278 ;
  assign n25281 = n25279 | n25280 ;
  assign n25282 = n25274 | n25281 ;
  assign n25283 = n25274 & n25281 ;
  assign n33668 = ~n25283 ;
  assign n25284 = n25282 & n33668 ;
  assign n33669 = ~n25138 ;
  assign n25285 = n25100 & n33669 ;
  assign n25286 = n25137 | n25285 ;
  assign n25287 = n25284 | n25286 ;
  assign n25288 = n25284 & n25286 ;
  assign n33670 = ~n25288 ;
  assign n25289 = n25287 & n33670 ;
  assign n4451 = n1690 & n4442 ;
  assign n1581 = x[110] & n1551 ;
  assign n1625 = x[111] & n1616 ;
  assign n25290 = n1581 | n1625 ;
  assign n25291 = x[112] & n1547 ;
  assign n25292 = n25290 | n25291 ;
  assign n25293 = n4451 | n25292 ;
  assign n33671 = ~n25293 ;
  assign n25294 = x[53] & n33671 ;
  assign n25295 = n30125 & n25293 ;
  assign n25296 = n25294 | n25295 ;
  assign n25297 = n25289 | n25296 ;
  assign n25298 = n25289 & n25296 ;
  assign n33672 = ~n25298 ;
  assign n25299 = n25297 & n33672 ;
  assign n33673 = ~n25141 ;
  assign n25300 = n25093 & n33673 ;
  assign n33674 = ~n25144 ;
  assign n25301 = n33674 & n25151 ;
  assign n25302 = n25300 | n25301 ;
  assign n25303 = n25299 | n25302 ;
  assign n25304 = n25299 & n25302 ;
  assign n33675 = ~n25304 ;
  assign n25305 = n25303 & n33675 ;
  assign n4483 = n2007 & n4474 ;
  assign n1906 = x[113] & n1866 ;
  assign n1979 = x[114] & n1931 ;
  assign n25306 = n1906 | n1979 ;
  assign n25307 = x[115] & n1862 ;
  assign n25308 = n25306 | n25307 ;
  assign n25309 = n4483 | n25308 ;
  assign n33676 = ~n25309 ;
  assign n25310 = x[50] & n33676 ;
  assign n25311 = n29865 & n25309 ;
  assign n25312 = n25310 | n25311 ;
  assign n25313 = n25305 | n25312 ;
  assign n25314 = n25305 & n25312 ;
  assign n33677 = ~n25314 ;
  assign n25315 = n25313 & n33677 ;
  assign n33678 = ~n25315 ;
  assign n25316 = n25240 & n33678 ;
  assign n33679 = ~n25240 ;
  assign n25317 = n33679 & n25315 ;
  assign n25318 = n25316 | n25317 ;
  assign n33680 = ~n25318 ;
  assign n25319 = n25238 & n33680 ;
  assign n33681 = ~n25238 ;
  assign n25320 = n33681 & n25318 ;
  assign n25321 = n25319 | n25320 ;
  assign n33682 = ~n25321 ;
  assign n25322 = n25231 & n33682 ;
  assign n33683 = ~n25231 ;
  assign n25323 = n33683 & n25321 ;
  assign n25324 = n25322 | n25323 ;
  assign n4994 = n2635 & n4985 ;
  assign n2494 = x[119] & n2492 ;
  assign n2603 = x[120] & n2557 ;
  assign n25325 = n2494 | n2603 ;
  assign n25326 = x[121] & n2488 ;
  assign n25327 = n25325 | n25326 ;
  assign n25328 = n4994 | n25327 ;
  assign n33684 = ~n25328 ;
  assign n25329 = x[44] & n33684 ;
  assign n25330 = n29400 & n25328 ;
  assign n25331 = n25329 | n25330 ;
  assign n25332 = n25324 | n25331 ;
  assign n25333 = n25324 & n25331 ;
  assign n33685 = ~n25333 ;
  assign n25334 = n25332 & n33685 ;
  assign n33686 = ~n25187 ;
  assign n25335 = n25087 & n33686 ;
  assign n25336 = n25186 | n25335 ;
  assign n25337 = n25334 | n25336 ;
  assign n25338 = n25334 & n25336 ;
  assign n33687 = ~n25338 ;
  assign n25339 = n25337 & n33687 ;
  assign n5845 = n3162 & n5838 ;
  assign n3032 = x[122] & n3031 ;
  assign n3137 = x[123] & n3096 ;
  assign n25340 = n3032 | n3137 ;
  assign n25341 = x[124] & n3027 ;
  assign n25342 = n25340 | n25341 ;
  assign n25343 = n5845 | n25342 ;
  assign n33688 = ~n25343 ;
  assign n25344 = x[41] & n33688 ;
  assign n25345 = n29184 & n25343 ;
  assign n25346 = n25344 | n25345 ;
  assign n25347 = n25339 | n25346 ;
  assign n25348 = n25339 & n25346 ;
  assign n33689 = ~n25348 ;
  assign n25349 = n25347 & n33689 ;
  assign n33690 = ~n25193 ;
  assign n25350 = n33690 & n25200 ;
  assign n25351 = n25191 | n25350 ;
  assign n33691 = ~n25351 ;
  assign n25352 = n25349 & n33691 ;
  assign n33692 = ~n25349 ;
  assign n25353 = n33692 & n25351 ;
  assign n25354 = n25352 | n25353 ;
  assign n5637 = n3574 & n5629 ;
  assign n3473 = x[125] & n3443 ;
  assign n3514 = x[126] & n3508 ;
  assign n25355 = n3473 | n3514 ;
  assign n25356 = x[127] & n3439 ;
  assign n25357 = n25355 | n25356 ;
  assign n25358 = n5637 | n25357 ;
  assign n33693 = ~n25358 ;
  assign n25359 = x[38] & n33693 ;
  assign n25360 = n28996 & n25358 ;
  assign n25361 = n25359 | n25360 ;
  assign n25362 = n25354 | n25361 ;
  assign n25363 = n25354 & n25361 ;
  assign n33694 = ~n25363 ;
  assign n25364 = n25362 & n33694 ;
  assign n33695 = ~n25208 ;
  assign n25365 = n33695 & n25215 ;
  assign n25366 = n25207 | n25365 ;
  assign n25367 = n25364 | n25366 ;
  assign n25368 = n25364 & n25366 ;
  assign n33696 = ~n25368 ;
  assign n25369 = n25367 & n33696 ;
  assign n33697 = ~n25218 ;
  assign n25219 = n25078 & n33697 ;
  assign n25370 = n25077 | n25219 ;
  assign n25371 = n25369 | n25370 ;
  assign n25372 = n25369 & n25370 ;
  assign n33698 = ~n25372 ;
  assign n25373 = n25371 & n33698 ;
  assign n25374 = n25229 & n25373 ;
  assign n25375 = n25229 | n25373 ;
  assign n33699 = ~n25374 ;
  assign n228 = n33699 & n25375 ;
  assign n33700 = ~n25339 ;
  assign n25499 = n33700 & n25346 ;
  assign n25500 = n25353 | n25499 ;
  assign n6188 = n3574 & n6186 ;
  assign n3507 = x[126] & n3443 ;
  assign n25501 = x[127] & n3508 ;
  assign n25502 = n3507 | n25501 ;
  assign n25503 = n6188 | n25502 ;
  assign n33701 = ~n25503 ;
  assign n25504 = x[38] & n33701 ;
  assign n25505 = n28996 & n25503 ;
  assign n25506 = n25504 | n25505 ;
  assign n25507 = n25500 | n25506 ;
  assign n25508 = n25500 & n25506 ;
  assign n33702 = ~n25508 ;
  assign n25509 = n25507 & n33702 ;
  assign n3008 = n1006 & n3001 ;
  assign n937 = x[102] & n900 ;
  assign n952 = x[103] & n949 ;
  assign n25377 = n937 | n952 ;
  assign n25378 = x[104] & n881 ;
  assign n25379 = n25377 | n25378 ;
  assign n25380 = n3008 | n25379 ;
  assign n33703 = ~n25380 ;
  assign n25381 = x[62] & n33703 ;
  assign n25382 = n30886 & n25380 ;
  assign n25383 = n25381 | n25382 ;
  assign n291 = x[100] & n27215 ;
  assign n821 = x[101] & n805 ;
  assign n25384 = n291 | n821 ;
  assign n25386 = n28822 & n25102 ;
  assign n25387 = n25245 | n25386 ;
  assign n25388 = n25384 | n25387 ;
  assign n25389 = n25384 & n25387 ;
  assign n33704 = ~n25389 ;
  assign n25390 = n25388 & n33704 ;
  assign n33705 = ~n25383 ;
  assign n25391 = n33705 & n25390 ;
  assign n33706 = ~n25390 ;
  assign n25392 = n25383 & n33706 ;
  assign n25393 = n25391 | n25392 ;
  assign n33707 = ~n25249 ;
  assign n25394 = n33707 & n25256 ;
  assign n25395 = n25247 | n25394 ;
  assign n25396 = n25393 | n25395 ;
  assign n25397 = n25393 & n25395 ;
  assign n33708 = ~n25397 ;
  assign n25398 = n25396 & n33708 ;
  assign n3208 = n1217 & n3199 ;
  assign n1092 = x[105] & n1079 ;
  assign n1156 = x[106] & n1144 ;
  assign n25399 = n1092 | n1156 ;
  assign n25400 = x[107] & n1075 ;
  assign n25401 = n25399 | n25400 ;
  assign n25402 = n3208 | n25401 ;
  assign n33709 = ~n25402 ;
  assign n25403 = x[59] & n33709 ;
  assign n25404 = n30638 & n25402 ;
  assign n25405 = n25403 | n25404 ;
  assign n25406 = n25398 | n25405 ;
  assign n25407 = n25398 & n25405 ;
  assign n33710 = ~n25407 ;
  assign n25408 = n25406 & n33710 ;
  assign n33711 = ~n25259 ;
  assign n25409 = n33711 & n25266 ;
  assign n25410 = n25273 | n25409 ;
  assign n33712 = ~n25410 ;
  assign n25411 = n25408 & n33712 ;
  assign n33713 = ~n25408 ;
  assign n25412 = n33713 & n25410 ;
  assign n25413 = n25411 | n25412 ;
  assign n3622 = n1457 & n3615 ;
  assign n1332 = x[108] & n1319 ;
  assign n1394 = x[109] & n1384 ;
  assign n25414 = n1332 | n1394 ;
  assign n25415 = x[110] & n1315 ;
  assign n25416 = n25414 | n25415 ;
  assign n25417 = n3622 | n25416 ;
  assign n33714 = ~n25417 ;
  assign n25418 = x[56] & n33714 ;
  assign n25419 = n30379 & n25417 ;
  assign n25420 = n25418 | n25419 ;
  assign n25421 = n25413 | n25420 ;
  assign n25422 = n25413 & n25420 ;
  assign n33715 = ~n25422 ;
  assign n25423 = n25421 & n33715 ;
  assign n33716 = ~n25274 ;
  assign n25424 = n33716 & n25281 ;
  assign n33717 = ~n25284 ;
  assign n25425 = n33717 & n25286 ;
  assign n25426 = n25424 | n25425 ;
  assign n33718 = ~n25426 ;
  assign n25427 = n25423 & n33718 ;
  assign n33719 = ~n25423 ;
  assign n25428 = n33719 & n25426 ;
  assign n25429 = n25427 | n25428 ;
  assign n4098 = n1690 & n4087 ;
  assign n1584 = x[111] & n1551 ;
  assign n1624 = x[112] & n1616 ;
  assign n25430 = n1584 | n1624 ;
  assign n25431 = x[113] & n1547 ;
  assign n25432 = n25430 | n25431 ;
  assign n25433 = n4098 | n25432 ;
  assign n33720 = ~n25433 ;
  assign n25434 = x[53] & n33720 ;
  assign n25435 = n30125 & n25433 ;
  assign n25436 = n25434 | n25435 ;
  assign n25437 = n25429 | n25436 ;
  assign n25438 = n25429 & n25436 ;
  assign n33721 = ~n25438 ;
  assign n25439 = n25437 & n33721 ;
  assign n33722 = ~n25289 ;
  assign n25440 = n33722 & n25296 ;
  assign n33723 = ~n25299 ;
  assign n25441 = n33723 & n25302 ;
  assign n25442 = n25440 | n25441 ;
  assign n33724 = ~n25442 ;
  assign n25443 = n25439 & n33724 ;
  assign n33725 = ~n25439 ;
  assign n25444 = n33725 & n25442 ;
  assign n25445 = n25443 | n25444 ;
  assign n4710 = n2007 & n4702 ;
  assign n1895 = x[114] & n1866 ;
  assign n1937 = x[115] & n1931 ;
  assign n25446 = n1895 | n1937 ;
  assign n25447 = x[116] & n1862 ;
  assign n25448 = n25446 | n25447 ;
  assign n25449 = n4710 | n25448 ;
  assign n33726 = ~n25449 ;
  assign n25450 = x[50] & n33726 ;
  assign n25451 = n29865 & n25449 ;
  assign n25452 = n25450 | n25451 ;
  assign n25453 = n25445 | n25452 ;
  assign n25454 = n25445 & n25452 ;
  assign n33727 = ~n25454 ;
  assign n25455 = n25453 & n33727 ;
  assign n33728 = ~n25305 ;
  assign n25456 = n33728 & n25312 ;
  assign n25457 = n25316 | n25456 ;
  assign n33729 = ~n25457 ;
  assign n25458 = n25455 & n33729 ;
  assign n33730 = ~n25455 ;
  assign n25459 = n33730 & n25457 ;
  assign n25460 = n25458 | n25459 ;
  assign n5057 = n2321 & n5047 ;
  assign n2232 = x[117] & n2179 ;
  assign n2246 = x[118] & n2244 ;
  assign n25461 = n2232 | n2246 ;
  assign n25462 = x[119] & n2175 ;
  assign n25463 = n25461 | n25462 ;
  assign n25464 = n5057 | n25463 ;
  assign n33731 = ~n25464 ;
  assign n25465 = x[47] & n33731 ;
  assign n25466 = n29621 & n25464 ;
  assign n25467 = n25465 | n25466 ;
  assign n33732 = ~n25467 ;
  assign n25468 = n25460 & n33732 ;
  assign n33733 = ~n25460 ;
  assign n25469 = n33733 & n25467 ;
  assign n25470 = n25468 | n25469 ;
  assign n25471 = n25319 | n25322 ;
  assign n25472 = n25470 | n25471 ;
  assign n25473 = n25470 & n25471 ;
  assign n33734 = ~n25473 ;
  assign n25474 = n25472 & n33734 ;
  assign n5025 = n2635 & n5022 ;
  assign n2527 = x[120] & n2492 ;
  assign n2559 = x[121] & n2557 ;
  assign n25475 = n2527 | n2559 ;
  assign n25476 = x[122] & n2488 ;
  assign n25477 = n25475 | n25476 ;
  assign n25478 = n5025 | n25477 ;
  assign n33735 = ~n25478 ;
  assign n25479 = x[44] & n33735 ;
  assign n25480 = n29400 & n25478 ;
  assign n25481 = n25479 | n25480 ;
  assign n25482 = n25474 | n25481 ;
  assign n25483 = n25474 & n25481 ;
  assign n33736 = ~n25483 ;
  assign n25484 = n25482 & n33736 ;
  assign n33737 = ~n25324 ;
  assign n25485 = n33737 & n25331 ;
  assign n33738 = ~n25334 ;
  assign n25486 = n33738 & n25336 ;
  assign n25487 = n25485 | n25486 ;
  assign n33739 = ~n25487 ;
  assign n25488 = n25484 & n33739 ;
  assign n33740 = ~n25484 ;
  assign n25489 = n33740 & n25487 ;
  assign n25490 = n25488 | n25489 ;
  assign n3195 = n642 & n3162 ;
  assign n3087 = x[123] & n3031 ;
  assign n3157 = x[124] & n3096 ;
  assign n25491 = n3087 | n3157 ;
  assign n25492 = x[125] & n3027 ;
  assign n25493 = n25491 | n25492 ;
  assign n25494 = n3195 | n25493 ;
  assign n33741 = ~n25494 ;
  assign n25495 = x[41] & n33741 ;
  assign n25496 = n29184 & n25494 ;
  assign n25497 = n25495 | n25496 ;
  assign n33742 = ~n25490 ;
  assign n25498 = n33742 & n25497 ;
  assign n33743 = ~n25497 ;
  assign n25510 = n25490 & n33743 ;
  assign n33744 = ~n25510 ;
  assign n25511 = n25509 & n33744 ;
  assign n33745 = ~n25498 ;
  assign n25512 = n33745 & n25511 ;
  assign n33746 = ~n25512 ;
  assign n25513 = n25509 & n33746 ;
  assign n25514 = n25510 | n25512 ;
  assign n25515 = n25498 | n25514 ;
  assign n33747 = ~n25513 ;
  assign n25516 = n33747 & n25515 ;
  assign n33748 = ~n25354 ;
  assign n25517 = n33748 & n25361 ;
  assign n33749 = ~n25364 ;
  assign n25518 = n33749 & n25366 ;
  assign n25519 = n25517 | n25518 ;
  assign n33750 = ~n25519 ;
  assign n25520 = n25516 & n33750 ;
  assign n33751 = ~n25516 ;
  assign n25521 = n33751 & n25519 ;
  assign n25522 = n25520 | n25521 ;
  assign n33752 = ~n25369 ;
  assign n25523 = n33752 & n25370 ;
  assign n33753 = ~n25523 ;
  assign n25524 = n25375 & n33753 ;
  assign n25525 = n25522 | n25524 ;
  assign n25526 = n25522 & n25524 ;
  assign n33754 = ~n25526 ;
  assign n229 = n25525 & n33754 ;
  assign n33755 = ~n25521 ;
  assign n25528 = n33755 & n25525 ;
  assign n25529 = n25508 | n25512 ;
  assign n25530 = n25489 | n25498 ;
  assign n3498 = x[127] & n3443 ;
  assign n5362 = n3574 & n5360 ;
  assign n25531 = n3498 | n5362 ;
  assign n33756 = ~n25531 ;
  assign n25532 = x[38] & n33756 ;
  assign n25533 = n28996 & n25531 ;
  assign n25534 = n25532 | n25533 ;
  assign n25535 = n25530 | n25534 ;
  assign n25536 = n25530 & n25534 ;
  assign n33757 = ~n25536 ;
  assign n25537 = n25535 & n33757 ;
  assign n25538 = n25459 | n25469 ;
  assign n4687 = n2321 & n4678 ;
  assign n2223 = x[118] & n2179 ;
  assign n2287 = x[119] & n2244 ;
  assign n25539 = n2223 | n2287 ;
  assign n25540 = x[120] & n2175 ;
  assign n25541 = n25539 | n25540 ;
  assign n25542 = n4687 | n25541 ;
  assign n33758 = ~n25542 ;
  assign n25543 = x[47] & n33758 ;
  assign n25544 = n29621 & n25542 ;
  assign n25545 = n25543 | n25544 ;
  assign n33759 = ~n25445 ;
  assign n25546 = n33759 & n25452 ;
  assign n25547 = n25444 | n25546 ;
  assign n2021 = n797 & n2007 ;
  assign n1873 = x[115] & n1866 ;
  assign n1936 = x[116] & n1931 ;
  assign n25612 = n1873 | n1936 ;
  assign n25613 = x[117] & n1862 ;
  assign n25614 = n25612 | n25613 ;
  assign n25615 = n2021 | n25614 ;
  assign n25616 = x[50] | n25615 ;
  assign n25617 = x[50] & n25615 ;
  assign n33760 = ~n25617 ;
  assign n25618 = n25616 & n33760 ;
  assign n33761 = ~n25429 ;
  assign n25548 = n33761 & n25436 ;
  assign n25549 = n25428 | n25548 ;
  assign n33762 = ~n25384 ;
  assign n25550 = n33762 & n25387 ;
  assign n25551 = n25392 | n25550 ;
  assign n292 = x[101] & n27215 ;
  assign n820 = x[102] & n805 ;
  assign n25552 = n292 | n820 ;
  assign n25553 = n25384 | n25552 ;
  assign n25554 = n25384 & n25552 ;
  assign n33763 = ~n25554 ;
  assign n25555 = n25553 & n33763 ;
  assign n33764 = ~n25551 ;
  assign n25556 = n33764 & n25555 ;
  assign n33765 = ~n25555 ;
  assign n25557 = n25551 & n33765 ;
  assign n25558 = n25556 | n25557 ;
  assign n3419 = n1006 & n3409 ;
  assign n939 = x[103] & n900 ;
  assign n960 = x[104] & n949 ;
  assign n25559 = n939 | n960 ;
  assign n25560 = x[105] & n881 ;
  assign n25561 = n25559 | n25560 ;
  assign n25562 = n3419 | n25561 ;
  assign n33766 = ~n25562 ;
  assign n25563 = x[62] & n33766 ;
  assign n25564 = n30886 & n25562 ;
  assign n25565 = n25563 | n25564 ;
  assign n33767 = ~n25565 ;
  assign n25566 = n25558 & n33767 ;
  assign n33768 = ~n25558 ;
  assign n25567 = n33768 & n25565 ;
  assign n25568 = n25566 | n25567 ;
  assign n3884 = n1217 & n3876 ;
  assign n1091 = x[106] & n1079 ;
  assign n1172 = x[107] & n1144 ;
  assign n25569 = n1091 | n1172 ;
  assign n25570 = x[108] & n1075 ;
  assign n25571 = n25569 | n25570 ;
  assign n25572 = n3884 | n25571 ;
  assign n33769 = ~n25572 ;
  assign n25573 = x[59] & n33769 ;
  assign n25574 = n30638 & n25572 ;
  assign n25575 = n25573 | n25574 ;
  assign n33770 = ~n25575 ;
  assign n25576 = n25568 & n33770 ;
  assign n33771 = ~n25568 ;
  assign n25577 = n33771 & n25575 ;
  assign n25578 = n25576 | n25577 ;
  assign n33772 = ~n25393 ;
  assign n25579 = n33772 & n25395 ;
  assign n33773 = ~n25398 ;
  assign n25580 = n33773 & n25405 ;
  assign n25581 = n25579 | n25580 ;
  assign n33774 = ~n25581 ;
  assign n25582 = n25578 & n33774 ;
  assign n33775 = ~n25578 ;
  assign n25583 = n33775 & n25581 ;
  assign n25584 = n25582 | n25583 ;
  assign n4250 = n1457 & n4246 ;
  assign n1331 = x[109] & n1319 ;
  assign n1393 = x[110] & n1384 ;
  assign n25585 = n1331 | n1393 ;
  assign n25586 = x[111] & n1315 ;
  assign n25587 = n25585 | n25586 ;
  assign n25588 = n4250 | n25587 ;
  assign n33776 = ~n25588 ;
  assign n25589 = x[56] & n33776 ;
  assign n25590 = n30379 & n25588 ;
  assign n25591 = n25589 | n25590 ;
  assign n25592 = n25584 | n25591 ;
  assign n25593 = n25584 & n25591 ;
  assign n33777 = ~n25593 ;
  assign n25594 = n25592 & n33777 ;
  assign n33778 = ~n25413 ;
  assign n25595 = n33778 & n25420 ;
  assign n25596 = n25412 | n25595 ;
  assign n33779 = ~n25596 ;
  assign n25597 = n25594 & n33779 ;
  assign n33780 = ~n25594 ;
  assign n25598 = n33780 & n25596 ;
  assign n25599 = n25597 | n25598 ;
  assign n4285 = n1690 & n4276 ;
  assign n1572 = x[112] & n1551 ;
  assign n1651 = x[113] & n1616 ;
  assign n25600 = n1572 | n1651 ;
  assign n25601 = x[114] & n1547 ;
  assign n25602 = n25600 | n25601 ;
  assign n25603 = n4285 | n25602 ;
  assign n33781 = ~n25603 ;
  assign n25604 = x[53] & n33781 ;
  assign n25605 = n30125 & n25603 ;
  assign n25606 = n25604 | n25605 ;
  assign n25607 = n25599 | n25606 ;
  assign n25608 = n25599 & n25606 ;
  assign n33782 = ~n25608 ;
  assign n25609 = n25607 & n33782 ;
  assign n25610 = n25549 | n25609 ;
  assign n25611 = n25549 & n25609 ;
  assign n33783 = ~n25611 ;
  assign n25619 = n25610 & n33783 ;
  assign n33784 = ~n25619 ;
  assign n25620 = n25618 & n33784 ;
  assign n33785 = ~n25618 ;
  assign n25621 = n25610 & n33785 ;
  assign n25622 = n33783 & n25621 ;
  assign n25623 = n25620 | n25622 ;
  assign n33786 = ~n25547 ;
  assign n25624 = n33786 & n25623 ;
  assign n33787 = ~n25623 ;
  assign n25625 = n25547 & n33787 ;
  assign n25626 = n25624 | n25625 ;
  assign n25627 = n25545 | n25626 ;
  assign n25628 = n25545 & n25626 ;
  assign n33788 = ~n25628 ;
  assign n25629 = n25627 & n33788 ;
  assign n25630 = n25538 | n25629 ;
  assign n25631 = n25538 & n25629 ;
  assign n33789 = ~n25631 ;
  assign n25632 = n25630 & n33789 ;
  assign n5422 = n2635 & n5417 ;
  assign n2493 = x[121] & n2492 ;
  assign n2615 = x[122] & n2557 ;
  assign n25633 = n2493 | n2615 ;
  assign n25634 = x[123] & n2488 ;
  assign n25635 = n25633 | n25634 ;
  assign n25636 = n5422 | n25635 ;
  assign n33790 = ~n25636 ;
  assign n25637 = x[44] & n33790 ;
  assign n25638 = n29400 & n25636 ;
  assign n25639 = n25637 | n25638 ;
  assign n25640 = n25632 | n25639 ;
  assign n25641 = n25632 & n25639 ;
  assign n33791 = ~n25641 ;
  assign n25642 = n25640 & n33791 ;
  assign n33792 = ~n25470 ;
  assign n25643 = n33792 & n25471 ;
  assign n33793 = ~n25474 ;
  assign n25644 = n33793 & n25481 ;
  assign n25645 = n25643 | n25644 ;
  assign n33794 = ~n25645 ;
  assign n25646 = n25642 & n33794 ;
  assign n33795 = ~n25642 ;
  assign n25647 = n33795 & n25645 ;
  assign n25648 = n25646 | n25647 ;
  assign n5390 = n3162 & n5388 ;
  assign n3093 = x[124] & n3031 ;
  assign n3158 = x[125] & n3096 ;
  assign n25649 = n3093 | n3158 ;
  assign n25650 = x[126] & n3027 ;
  assign n25651 = n25649 | n25650 ;
  assign n25652 = n5390 | n25651 ;
  assign n33796 = ~n25652 ;
  assign n25653 = x[41] & n33796 ;
  assign n25654 = n29184 & n25652 ;
  assign n25655 = n25653 | n25654 ;
  assign n25656 = n25648 | n25655 ;
  assign n25657 = n25648 & n25655 ;
  assign n33797 = ~n25657 ;
  assign n25658 = n25656 & n33797 ;
  assign n25660 = n25537 & n25658 ;
  assign n25661 = n25537 | n25658 ;
  assign n33798 = ~n25660 ;
  assign n25662 = n33798 & n25661 ;
  assign n33799 = ~n25529 ;
  assign n25663 = n33799 & n25662 ;
  assign n33800 = ~n25662 ;
  assign n25664 = n25529 & n33800 ;
  assign n25665 = n25663 | n25664 ;
  assign n25666 = n25528 & n25665 ;
  assign n25667 = n25528 | n25665 ;
  assign n33801 = ~n25666 ;
  assign n230 = n33801 & n25667 ;
  assign n33802 = ~n25664 ;
  assign n25669 = n33802 & n25667 ;
  assign n33803 = ~n25609 ;
  assign n25670 = n25549 & n33803 ;
  assign n25671 = n25620 | n25670 ;
  assign n2008 = n784 & n2007 ;
  assign n1871 = x[116] & n1866 ;
  assign n1984 = x[117] & n1931 ;
  assign n25672 = n1871 | n1984 ;
  assign n25673 = x[118] & n1862 ;
  assign n25674 = n25672 | n25673 ;
  assign n25675 = n2008 | n25674 ;
  assign n25676 = x[50] | n25675 ;
  assign n25677 = x[50] & n25675 ;
  assign n33804 = ~n25677 ;
  assign n25678 = n25676 & n33804 ;
  assign n33805 = ~n25599 ;
  assign n25679 = n33805 & n25606 ;
  assign n25680 = n25598 | n25679 ;
  assign n25681 = n33762 & n25552 ;
  assign n25682 = n25557 | n25681 ;
  assign n293 = x[102] & n27215 ;
  assign n818 = x[103] & n805 ;
  assign n25683 = n293 | n818 ;
  assign n25385 = x[38] | n25384 ;
  assign n25684 = x[38] & n25384 ;
  assign n33806 = ~n25684 ;
  assign n25685 = n25385 & n33806 ;
  assign n33807 = ~n25683 ;
  assign n25686 = n33807 & n25685 ;
  assign n33808 = ~n25685 ;
  assign n25687 = n25683 & n33808 ;
  assign n25688 = n25686 | n25687 ;
  assign n25689 = n25682 | n25688 ;
  assign n25690 = n25682 & n25688 ;
  assign n33809 = ~n25690 ;
  assign n25691 = n25689 & n33809 ;
  assign n3224 = n1006 & n3223 ;
  assign n940 = x[104] & n900 ;
  assign n971 = x[105] & n949 ;
  assign n25692 = n940 | n971 ;
  assign n25693 = x[106] & n881 ;
  assign n25694 = n25692 | n25693 ;
  assign n25695 = n3224 | n25694 ;
  assign n33810 = ~n25695 ;
  assign n25696 = x[62] & n33810 ;
  assign n25697 = n30886 & n25695 ;
  assign n25698 = n25696 | n25697 ;
  assign n25699 = n25691 | n25698 ;
  assign n25700 = n25691 & n25698 ;
  assign n33811 = ~n25700 ;
  assign n25701 = n25699 & n33811 ;
  assign n3649 = n1217 & n3639 ;
  assign n1090 = x[107] & n1079 ;
  assign n1154 = x[108] & n1144 ;
  assign n25702 = n1090 | n1154 ;
  assign n25703 = x[109] & n1075 ;
  assign n25704 = n25702 | n25703 ;
  assign n25705 = n3649 | n25704 ;
  assign n33812 = ~n25705 ;
  assign n25706 = x[59] & n33812 ;
  assign n25707 = n30638 & n25705 ;
  assign n25708 = n25706 | n25707 ;
  assign n33813 = ~n25708 ;
  assign n25709 = n25701 & n33813 ;
  assign n33814 = ~n25701 ;
  assign n25710 = n33814 & n25708 ;
  assign n25711 = n25709 | n25710 ;
  assign n25712 = n25567 | n25577 ;
  assign n25713 = n25711 | n25712 ;
  assign n25714 = n25711 & n25712 ;
  assign n33815 = ~n25714 ;
  assign n25715 = n25713 & n33815 ;
  assign n4452 = n1457 & n4442 ;
  assign n1322 = x[110] & n1319 ;
  assign n1391 = x[111] & n1384 ;
  assign n25716 = n1322 | n1391 ;
  assign n25717 = x[112] & n1315 ;
  assign n25718 = n25716 | n25717 ;
  assign n25719 = n4452 | n25718 ;
  assign n33816 = ~n25719 ;
  assign n25720 = x[56] & n33816 ;
  assign n25721 = n30379 & n25719 ;
  assign n25722 = n25720 | n25721 ;
  assign n25723 = n25715 | n25722 ;
  assign n25724 = n25715 & n25722 ;
  assign n33817 = ~n25724 ;
  assign n25725 = n25723 & n33817 ;
  assign n33818 = ~n25584 ;
  assign n25726 = n33818 & n25591 ;
  assign n25727 = n25583 | n25726 ;
  assign n25728 = n25725 | n25727 ;
  assign n25729 = n25725 & n25727 ;
  assign n33819 = ~n25729 ;
  assign n25730 = n25728 & n33819 ;
  assign n4484 = n1690 & n4474 ;
  assign n1559 = x[113] & n1551 ;
  assign n1627 = x[114] & n1616 ;
  assign n25731 = n1559 | n1627 ;
  assign n25732 = x[115] & n1547 ;
  assign n25733 = n25731 | n25732 ;
  assign n25734 = n4484 | n25733 ;
  assign n33820 = ~n25734 ;
  assign n25735 = x[53] & n33820 ;
  assign n25736 = n30125 & n25734 ;
  assign n25737 = n25735 | n25736 ;
  assign n25738 = n25730 | n25737 ;
  assign n25739 = n25730 & n25737 ;
  assign n33821 = ~n25739 ;
  assign n25740 = n25738 & n33821 ;
  assign n33822 = ~n25740 ;
  assign n25741 = n25680 & n33822 ;
  assign n33823 = ~n25680 ;
  assign n25742 = n33823 & n25740 ;
  assign n25743 = n25741 | n25742 ;
  assign n33824 = ~n25743 ;
  assign n25744 = n25678 & n33824 ;
  assign n33825 = ~n25678 ;
  assign n25745 = n33825 & n25743 ;
  assign n25746 = n25744 | n25745 ;
  assign n33826 = ~n25746 ;
  assign n25747 = n25671 & n33826 ;
  assign n33827 = ~n25671 ;
  assign n25748 = n33827 & n25746 ;
  assign n25749 = n25747 | n25748 ;
  assign n4989 = n2321 & n4985 ;
  assign n2180 = x[119] & n2179 ;
  assign n2294 = x[120] & n2244 ;
  assign n25750 = n2180 | n2294 ;
  assign n25751 = x[121] & n2175 ;
  assign n25752 = n25750 | n25751 ;
  assign n25753 = n4989 | n25752 ;
  assign n33828 = ~n25753 ;
  assign n25754 = x[47] & n33828 ;
  assign n25755 = n29621 & n25753 ;
  assign n25756 = n25754 | n25755 ;
  assign n25757 = n25749 | n25756 ;
  assign n25758 = n25749 & n25756 ;
  assign n33829 = ~n25758 ;
  assign n25759 = n25757 & n33829 ;
  assign n33830 = ~n25626 ;
  assign n25760 = n25545 & n33830 ;
  assign n25761 = n25625 | n25760 ;
  assign n25762 = n25759 | n25761 ;
  assign n25763 = n25759 & n25761 ;
  assign n33831 = ~n25763 ;
  assign n25764 = n25762 & n33831 ;
  assign n5840 = n2635 & n5838 ;
  assign n2518 = x[122] & n2492 ;
  assign n2558 = x[123] & n2557 ;
  assign n25765 = n2518 | n2558 ;
  assign n25766 = x[124] & n2488 ;
  assign n25767 = n25765 | n25766 ;
  assign n25768 = n5840 | n25767 ;
  assign n33832 = ~n25768 ;
  assign n25769 = x[44] & n33832 ;
  assign n25770 = n29400 & n25768 ;
  assign n25771 = n25769 | n25770 ;
  assign n25772 = n25764 | n25771 ;
  assign n25773 = n25764 & n25771 ;
  assign n33833 = ~n25773 ;
  assign n25774 = n25772 & n33833 ;
  assign n33834 = ~n25629 ;
  assign n25775 = n25538 & n33834 ;
  assign n33835 = ~n25632 ;
  assign n25776 = n33835 & n25639 ;
  assign n25777 = n25775 | n25776 ;
  assign n33836 = ~n25777 ;
  assign n25778 = n25774 & n33836 ;
  assign n33837 = ~n25774 ;
  assign n25779 = n33837 & n25777 ;
  assign n25780 = n25778 | n25779 ;
  assign n5642 = n3162 & n5629 ;
  assign n3094 = x[125] & n3031 ;
  assign n3111 = x[126] & n3096 ;
  assign n25781 = n3094 | n3111 ;
  assign n25782 = x[127] & n3027 ;
  assign n25783 = n25781 | n25782 ;
  assign n25784 = n5642 | n25783 ;
  assign n33838 = ~n25784 ;
  assign n25785 = x[41] & n33838 ;
  assign n25786 = n29184 & n25784 ;
  assign n25787 = n25785 | n25786 ;
  assign n25788 = n25780 | n25787 ;
  assign n25789 = n25780 & n25787 ;
  assign n33839 = ~n25789 ;
  assign n25790 = n25788 & n33839 ;
  assign n33840 = ~n25648 ;
  assign n25791 = n33840 & n25655 ;
  assign n25792 = n25647 | n25791 ;
  assign n25793 = n25790 | n25792 ;
  assign n25794 = n25790 & n25792 ;
  assign n33841 = ~n25794 ;
  assign n25795 = n25793 & n33841 ;
  assign n33842 = ~n25658 ;
  assign n25659 = n25537 & n33842 ;
  assign n25796 = n25536 | n25659 ;
  assign n25797 = n25795 | n25796 ;
  assign n25798 = n25795 & n25796 ;
  assign n33843 = ~n25798 ;
  assign n25799 = n25797 & n33843 ;
  assign n25800 = n25669 | n25799 ;
  assign n25801 = n25669 & n25799 ;
  assign n33844 = ~n25801 ;
  assign n231 = n25800 & n33844 ;
  assign n33845 = ~n25764 ;
  assign n25912 = n33845 & n25771 ;
  assign n25913 = n25779 | n25912 ;
  assign n6196 = n3162 & n6186 ;
  assign n3095 = x[126] & n3031 ;
  assign n25914 = x[127] & n3096 ;
  assign n25915 = n3095 | n25914 ;
  assign n25916 = n6196 | n25915 ;
  assign n33846 = ~n25916 ;
  assign n25917 = x[41] & n33846 ;
  assign n25918 = n29184 & n25916 ;
  assign n25919 = n25917 | n25918 ;
  assign n25920 = n25913 | n25919 ;
  assign n25921 = n25913 & n25919 ;
  assign n33847 = ~n25921 ;
  assign n25922 = n25920 & n33847 ;
  assign n33848 = ~n25688 ;
  assign n25803 = n25682 & n33848 ;
  assign n33849 = ~n25691 ;
  assign n25804 = n33849 & n25698 ;
  assign n25805 = n25803 | n25804 ;
  assign n294 = x[103] & n27215 ;
  assign n808 = x[104] & n805 ;
  assign n25806 = n294 | n808 ;
  assign n25808 = n28996 & n25384 ;
  assign n25809 = n25687 | n25808 ;
  assign n25810 = n25806 | n25809 ;
  assign n25811 = n25806 & n25809 ;
  assign n33850 = ~n25811 ;
  assign n25812 = n25810 & n33850 ;
  assign n882 = x[107] & n881 ;
  assign n25813 = x[105] & n900 ;
  assign n25814 = x[106] & n949 ;
  assign n25815 = n25813 | n25814 ;
  assign n25816 = n882 | n25815 ;
  assign n25817 = n1006 & n3199 ;
  assign n25818 = n25816 | n25817 ;
  assign n25819 = n30886 & n25818 ;
  assign n33851 = ~n25818 ;
  assign n25820 = x[62] & n33851 ;
  assign n25821 = n25819 | n25820 ;
  assign n25822 = n25812 | n25821 ;
  assign n25823 = n25812 & n25821 ;
  assign n33852 = ~n25823 ;
  assign n25824 = n25822 & n33852 ;
  assign n25825 = n25805 | n25824 ;
  assign n25826 = n25805 & n25824 ;
  assign n33853 = ~n25826 ;
  assign n25827 = n25825 & n33853 ;
  assign n3623 = n1217 & n3615 ;
  assign n1137 = x[108] & n1079 ;
  assign n1183 = x[109] & n1144 ;
  assign n25828 = n1137 | n1183 ;
  assign n25829 = x[110] & n1075 ;
  assign n25830 = n25828 | n25829 ;
  assign n25831 = n3623 | n25830 ;
  assign n33854 = ~n25831 ;
  assign n25832 = x[59] & n33854 ;
  assign n25833 = n30638 & n25831 ;
  assign n25834 = n25832 | n25833 ;
  assign n25835 = n25827 | n25834 ;
  assign n25836 = n25827 & n25834 ;
  assign n33855 = ~n25836 ;
  assign n25837 = n25835 & n33855 ;
  assign n33856 = ~n25711 ;
  assign n25838 = n33856 & n25712 ;
  assign n25839 = n25710 | n25838 ;
  assign n33857 = ~n25839 ;
  assign n25840 = n25837 & n33857 ;
  assign n33858 = ~n25837 ;
  assign n25841 = n33858 & n25839 ;
  assign n25842 = n25840 | n25841 ;
  assign n4099 = n1457 & n4087 ;
  assign n1327 = x[111] & n1319 ;
  assign n1442 = x[112] & n1384 ;
  assign n25843 = n1327 | n1442 ;
  assign n25844 = x[113] & n1315 ;
  assign n25845 = n25843 | n25844 ;
  assign n25846 = n4099 | n25845 ;
  assign n33859 = ~n25846 ;
  assign n25847 = x[56] & n33859 ;
  assign n25848 = n30379 & n25846 ;
  assign n25849 = n25847 | n25848 ;
  assign n25850 = n25842 | n25849 ;
  assign n25851 = n25842 & n25849 ;
  assign n33860 = ~n25851 ;
  assign n25852 = n25850 & n33860 ;
  assign n33861 = ~n25715 ;
  assign n25853 = n33861 & n25722 ;
  assign n33862 = ~n25725 ;
  assign n25854 = n33862 & n25727 ;
  assign n25855 = n25853 | n25854 ;
  assign n33863 = ~n25855 ;
  assign n25856 = n25852 & n33863 ;
  assign n33864 = ~n25852 ;
  assign n25857 = n33864 & n25855 ;
  assign n25858 = n25856 | n25857 ;
  assign n4712 = n1690 & n4702 ;
  assign n1558 = x[114] & n1551 ;
  assign n1622 = x[115] & n1616 ;
  assign n25859 = n1558 | n1622 ;
  assign n25860 = x[116] & n1547 ;
  assign n25861 = n25859 | n25860 ;
  assign n25862 = n4712 | n25861 ;
  assign n33865 = ~n25862 ;
  assign n25863 = x[53] & n33865 ;
  assign n25864 = n30125 & n25862 ;
  assign n25865 = n25863 | n25864 ;
  assign n25866 = n25858 | n25865 ;
  assign n25867 = n25858 & n25865 ;
  assign n33866 = ~n25867 ;
  assign n25868 = n25866 & n33866 ;
  assign n33867 = ~n25730 ;
  assign n25869 = n33867 & n25737 ;
  assign n25870 = n25741 | n25869 ;
  assign n33868 = ~n25870 ;
  assign n25871 = n25868 & n33868 ;
  assign n33869 = ~n25868 ;
  assign n25872 = n33869 & n25870 ;
  assign n25873 = n25871 | n25872 ;
  assign n5058 = n2007 & n5047 ;
  assign n1868 = x[117] & n1866 ;
  assign n1935 = x[118] & n1931 ;
  assign n25874 = n1868 | n1935 ;
  assign n25875 = x[119] & n1862 ;
  assign n25876 = n25874 | n25875 ;
  assign n25877 = n5058 | n25876 ;
  assign n33870 = ~n25877 ;
  assign n25878 = x[50] & n33870 ;
  assign n25879 = n29865 & n25877 ;
  assign n25880 = n25878 | n25879 ;
  assign n33871 = ~n25880 ;
  assign n25881 = n25873 & n33871 ;
  assign n33872 = ~n25873 ;
  assign n25882 = n33872 & n25880 ;
  assign n25883 = n25881 | n25882 ;
  assign n25884 = n25744 | n25747 ;
  assign n25885 = n25883 | n25884 ;
  assign n25886 = n25883 & n25884 ;
  assign n33873 = ~n25886 ;
  assign n25887 = n25885 & n33873 ;
  assign n5023 = n2321 & n5022 ;
  assign n2236 = x[120] & n2179 ;
  assign n2245 = x[121] & n2244 ;
  assign n25888 = n2236 | n2245 ;
  assign n25889 = x[122] & n2175 ;
  assign n25890 = n25888 | n25889 ;
  assign n25891 = n5023 | n25890 ;
  assign n33874 = ~n25891 ;
  assign n25892 = x[47] & n33874 ;
  assign n25893 = n29621 & n25891 ;
  assign n25894 = n25892 | n25893 ;
  assign n25895 = n25887 | n25894 ;
  assign n25896 = n25887 & n25894 ;
  assign n33875 = ~n25896 ;
  assign n25897 = n25895 & n33875 ;
  assign n33876 = ~n25749 ;
  assign n25898 = n33876 & n25756 ;
  assign n33877 = ~n25759 ;
  assign n25899 = n33877 & n25761 ;
  assign n25900 = n25898 | n25899 ;
  assign n33878 = ~n25900 ;
  assign n25901 = n25897 & n33878 ;
  assign n33879 = ~n25897 ;
  assign n25902 = n33879 & n25900 ;
  assign n25903 = n25901 | n25902 ;
  assign n2652 = n642 & n2635 ;
  assign n2555 = x[123] & n2492 ;
  assign n2617 = x[124] & n2557 ;
  assign n25904 = n2555 | n2617 ;
  assign n25905 = x[125] & n2488 ;
  assign n25906 = n25904 | n25905 ;
  assign n25907 = n2652 | n25906 ;
  assign n33880 = ~n25907 ;
  assign n25908 = x[44] & n33880 ;
  assign n25909 = n29400 & n25907 ;
  assign n25910 = n25908 | n25909 ;
  assign n33881 = ~n25903 ;
  assign n25911 = n33881 & n25910 ;
  assign n33882 = ~n25910 ;
  assign n25923 = n25903 & n33882 ;
  assign n33883 = ~n25923 ;
  assign n25924 = n25922 & n33883 ;
  assign n33884 = ~n25911 ;
  assign n25925 = n33884 & n25924 ;
  assign n33885 = ~n25925 ;
  assign n25926 = n25922 & n33885 ;
  assign n25927 = n25923 | n25925 ;
  assign n25928 = n25911 | n25927 ;
  assign n33886 = ~n25926 ;
  assign n25929 = n33886 & n25928 ;
  assign n33887 = ~n25780 ;
  assign n25930 = n33887 & n25787 ;
  assign n33888 = ~n25790 ;
  assign n25931 = n33888 & n25792 ;
  assign n25932 = n25930 | n25931 ;
  assign n33889 = ~n25932 ;
  assign n25933 = n25929 & n33889 ;
  assign n33890 = ~n25929 ;
  assign n25934 = n33890 & n25932 ;
  assign n25935 = n25933 | n25934 ;
  assign n33891 = ~n25795 ;
  assign n25936 = n33891 & n25796 ;
  assign n33892 = ~n25936 ;
  assign n25937 = n25800 & n33892 ;
  assign n25938 = n25935 & n25937 ;
  assign n25939 = n25935 | n25937 ;
  assign n33893 = ~n25938 ;
  assign n232 = n33893 & n25939 ;
  assign n33894 = ~n25934 ;
  assign n25941 = n33894 & n25939 ;
  assign n25942 = n25921 | n25925 ;
  assign n25943 = n25902 | n25911 ;
  assign n3082 = x[127] & n3031 ;
  assign n5369 = n3162 & n5360 ;
  assign n25944 = n3082 | n5369 ;
  assign n33895 = ~n25944 ;
  assign n25945 = x[41] & n33895 ;
  assign n25946 = n29184 & n25944 ;
  assign n25947 = n25945 | n25946 ;
  assign n25948 = n25943 | n25947 ;
  assign n25949 = n25943 & n25947 ;
  assign n33896 = ~n25949 ;
  assign n25950 = n25948 & n33896 ;
  assign n25951 = n25872 | n25882 ;
  assign n4688 = n2007 & n4678 ;
  assign n1921 = x[118] & n1866 ;
  assign n1981 = x[119] & n1931 ;
  assign n26017 = n1921 | n1981 ;
  assign n26018 = x[120] & n1862 ;
  assign n26019 = n26017 | n26018 ;
  assign n26020 = n4688 | n26019 ;
  assign n26021 = x[50] | n26020 ;
  assign n26022 = x[50] & n26020 ;
  assign n33897 = ~n26022 ;
  assign n26023 = n26021 & n33897 ;
  assign n33898 = ~n25858 ;
  assign n25952 = n33898 & n25865 ;
  assign n25953 = n25857 | n25952 ;
  assign n1695 = n797 & n1690 ;
  assign n1557 = x[115] & n1551 ;
  assign n1621 = x[116] & n1616 ;
  assign n26004 = n1557 | n1621 ;
  assign n26005 = x[117] & n1547 ;
  assign n26006 = n26004 | n26005 ;
  assign n26007 = n1695 | n26006 ;
  assign n26008 = x[53] | n26007 ;
  assign n26009 = x[53] & n26007 ;
  assign n33899 = ~n26009 ;
  assign n26010 = n26008 & n33899 ;
  assign n33900 = ~n25842 ;
  assign n25954 = n33900 & n25849 ;
  assign n25955 = n25841 | n25954 ;
  assign n33901 = ~n25824 ;
  assign n25956 = n25805 & n33901 ;
  assign n33902 = ~n25827 ;
  assign n25957 = n33902 & n25834 ;
  assign n25958 = n25956 | n25957 ;
  assign n33903 = ~n25806 ;
  assign n25959 = n33903 & n25809 ;
  assign n33904 = ~n25812 ;
  assign n25960 = n33904 & n25821 ;
  assign n25961 = n25959 | n25960 ;
  assign n295 = x[104] & n27215 ;
  assign n841 = x[105] & n805 ;
  assign n25962 = n295 | n841 ;
  assign n25963 = n25806 | n25962 ;
  assign n25964 = n25806 & n25962 ;
  assign n33905 = ~n25964 ;
  assign n25965 = n25963 & n33905 ;
  assign n33906 = ~n25961 ;
  assign n25966 = n33906 & n25965 ;
  assign n33907 = ~n25965 ;
  assign n25967 = n25961 & n33907 ;
  assign n25968 = n25966 | n25967 ;
  assign n3885 = n1006 & n3876 ;
  assign n928 = x[106] & n900 ;
  assign n973 = x[107] & n949 ;
  assign n25969 = n928 | n973 ;
  assign n25970 = x[108] & n881 ;
  assign n25971 = n25969 | n25970 ;
  assign n25972 = n3885 | n25971 ;
  assign n33908 = ~n25972 ;
  assign n25973 = x[62] & n33908 ;
  assign n25974 = n30886 & n25972 ;
  assign n25975 = n25973 | n25974 ;
  assign n33909 = ~n25975 ;
  assign n25976 = n25968 & n33909 ;
  assign n33910 = ~n25968 ;
  assign n25977 = n33910 & n25975 ;
  assign n25978 = n25976 | n25977 ;
  assign n4256 = n1217 & n4246 ;
  assign n1088 = x[109] & n1079 ;
  assign n1160 = x[110] & n1144 ;
  assign n25979 = n1088 | n1160 ;
  assign n25980 = x[111] & n1075 ;
  assign n25981 = n25979 | n25980 ;
  assign n25982 = n4256 | n25981 ;
  assign n33911 = ~n25982 ;
  assign n25983 = x[59] & n33911 ;
  assign n25984 = n30638 & n25982 ;
  assign n25985 = n25983 | n25984 ;
  assign n33912 = ~n25985 ;
  assign n25986 = n25978 & n33912 ;
  assign n33913 = ~n25978 ;
  assign n25987 = n33913 & n25985 ;
  assign n25988 = n25986 | n25987 ;
  assign n25989 = n25958 | n25988 ;
  assign n25990 = n25958 & n25988 ;
  assign n33914 = ~n25990 ;
  assign n25991 = n25989 & n33914 ;
  assign n4286 = n1457 & n4276 ;
  assign n1334 = x[112] & n1319 ;
  assign n1395 = x[113] & n1384 ;
  assign n25992 = n1334 | n1395 ;
  assign n25993 = x[114] & n1315 ;
  assign n25994 = n25992 | n25993 ;
  assign n25995 = n4286 | n25994 ;
  assign n33915 = ~n25995 ;
  assign n25996 = x[56] & n33915 ;
  assign n25997 = n30379 & n25995 ;
  assign n25998 = n25996 | n25997 ;
  assign n25999 = n25991 | n25998 ;
  assign n26000 = n25991 & n25998 ;
  assign n33916 = ~n26000 ;
  assign n26001 = n25999 & n33916 ;
  assign n26002 = n25955 | n26001 ;
  assign n26003 = n25955 & n26001 ;
  assign n33917 = ~n26003 ;
  assign n26011 = n26002 & n33917 ;
  assign n33918 = ~n26011 ;
  assign n26012 = n26010 & n33918 ;
  assign n33919 = ~n26010 ;
  assign n26013 = n26002 & n33919 ;
  assign n26014 = n33917 & n26013 ;
  assign n26015 = n26012 | n26014 ;
  assign n26016 = n25953 & n26015 ;
  assign n26024 = n25953 | n26015 ;
  assign n33920 = ~n26016 ;
  assign n26025 = n33920 & n26024 ;
  assign n33921 = ~n26025 ;
  assign n26026 = n26023 & n33921 ;
  assign n33922 = ~n26023 ;
  assign n26027 = n33922 & n26024 ;
  assign n26028 = n33920 & n26027 ;
  assign n26029 = n26026 | n26028 ;
  assign n33923 = ~n25951 ;
  assign n26030 = n33923 & n26029 ;
  assign n33924 = ~n26029 ;
  assign n26031 = n25951 & n33924 ;
  assign n26032 = n26030 | n26031 ;
  assign n5429 = n2321 & n5417 ;
  assign n2235 = x[121] & n2179 ;
  assign n2248 = x[122] & n2244 ;
  assign n26033 = n2235 | n2248 ;
  assign n26034 = x[123] & n2175 ;
  assign n26035 = n26033 | n26034 ;
  assign n26036 = n5429 | n26035 ;
  assign n33925 = ~n26036 ;
  assign n26037 = x[47] & n33925 ;
  assign n26038 = n29621 & n26036 ;
  assign n26039 = n26037 | n26038 ;
  assign n26040 = n26032 | n26039 ;
  assign n26041 = n26032 & n26039 ;
  assign n33926 = ~n26041 ;
  assign n26042 = n26040 & n33926 ;
  assign n33927 = ~n25883 ;
  assign n26043 = n33927 & n25884 ;
  assign n33928 = ~n25887 ;
  assign n26044 = n33928 & n25894 ;
  assign n26045 = n26043 | n26044 ;
  assign n33929 = ~n26045 ;
  assign n26046 = n26042 & n33929 ;
  assign n33930 = ~n26042 ;
  assign n26047 = n33930 & n26045 ;
  assign n26048 = n26046 | n26047 ;
  assign n5394 = n2635 & n5388 ;
  assign n2514 = x[124] & n2492 ;
  assign n2618 = x[125] & n2557 ;
  assign n26049 = n2514 | n2618 ;
  assign n26050 = x[126] & n2488 ;
  assign n26051 = n26049 | n26050 ;
  assign n26052 = n5394 | n26051 ;
  assign n33931 = ~n26052 ;
  assign n26053 = x[44] & n33931 ;
  assign n26054 = n29400 & n26052 ;
  assign n26055 = n26053 | n26054 ;
  assign n26056 = n26048 | n26055 ;
  assign n26057 = n26048 & n26055 ;
  assign n33932 = ~n26057 ;
  assign n26058 = n26056 & n33932 ;
  assign n26060 = n25950 & n26058 ;
  assign n26061 = n25950 | n26058 ;
  assign n33933 = ~n26060 ;
  assign n26062 = n33933 & n26061 ;
  assign n33934 = ~n25942 ;
  assign n26063 = n33934 & n26062 ;
  assign n33935 = ~n26062 ;
  assign n26064 = n25942 & n33935 ;
  assign n26065 = n26063 | n26064 ;
  assign n26066 = n25941 | n26065 ;
  assign n26067 = n25941 & n26065 ;
  assign n33936 = ~n26067 ;
  assign n233 = n26066 & n33936 ;
  assign n33937 = ~n26064 ;
  assign n26069 = n33937 & n26066 ;
  assign n33938 = ~n26015 ;
  assign n26070 = n25953 & n33938 ;
  assign n26071 = n26026 | n26070 ;
  assign n4996 = n2007 & n4985 ;
  assign n1880 = x[119] & n1866 ;
  assign n1962 = x[120] & n1931 ;
  assign n26072 = n1880 | n1962 ;
  assign n26073 = x[121] & n1862 ;
  assign n26074 = n26072 | n26073 ;
  assign n26075 = n4996 | n26074 ;
  assign n33939 = ~n26075 ;
  assign n26076 = x[50] & n33939 ;
  assign n26077 = n29865 & n26075 ;
  assign n26078 = n26076 | n26077 ;
  assign n33940 = ~n26001 ;
  assign n26079 = n25955 & n33940 ;
  assign n26080 = n26012 | n26079 ;
  assign n33941 = ~n25988 ;
  assign n26081 = n25958 & n33941 ;
  assign n33942 = ~n25991 ;
  assign n26082 = n33942 & n25998 ;
  assign n26083 = n26081 | n26082 ;
  assign n4476 = n1457 & n4474 ;
  assign n1329 = x[113] & n1319 ;
  assign n1389 = x[114] & n1384 ;
  assign n26084 = n1329 | n1389 ;
  assign n26085 = x[115] & n1315 ;
  assign n26086 = n26084 | n26085 ;
  assign n26087 = n4476 | n26086 ;
  assign n33943 = ~n26087 ;
  assign n26088 = x[56] & n33943 ;
  assign n26089 = n30379 & n26087 ;
  assign n26090 = n26088 | n26089 ;
  assign n25807 = x[41] | n25806 ;
  assign n26091 = x[41] & n25806 ;
  assign n33944 = ~n26091 ;
  assign n26092 = n25807 & n33944 ;
  assign n296 = x[105] & n27215 ;
  assign n838 = x[106] & n805 ;
  assign n26093 = n296 | n838 ;
  assign n33945 = ~n26093 ;
  assign n26094 = n26092 & n33945 ;
  assign n33946 = ~n26092 ;
  assign n26095 = n33946 & n26093 ;
  assign n26096 = n26094 | n26095 ;
  assign n3650 = n1006 & n3639 ;
  assign n941 = x[107] & n900 ;
  assign n990 = x[108] & n949 ;
  assign n26097 = n941 | n990 ;
  assign n26098 = x[109] & n881 ;
  assign n26099 = n26097 | n26098 ;
  assign n26100 = n3650 | n26099 ;
  assign n33947 = ~n26100 ;
  assign n26101 = x[62] & n33947 ;
  assign n26102 = n30886 & n26100 ;
  assign n26103 = n26101 | n26102 ;
  assign n26104 = n26096 | n26103 ;
  assign n26105 = n26096 & n26103 ;
  assign n33948 = ~n26105 ;
  assign n26106 = n26104 & n33948 ;
  assign n26107 = n33903 & n25962 ;
  assign n26108 = n25967 | n26107 ;
  assign n33949 = ~n26108 ;
  assign n26109 = n26106 & n33949 ;
  assign n33950 = ~n26106 ;
  assign n26110 = n33950 & n26108 ;
  assign n26111 = n26109 | n26110 ;
  assign n4453 = n1217 & n4442 ;
  assign n1087 = x[110] & n1079 ;
  assign n1191 = x[111] & n1144 ;
  assign n26112 = n1087 | n1191 ;
  assign n26113 = x[112] & n1075 ;
  assign n26114 = n26112 | n26113 ;
  assign n26115 = n4453 | n26114 ;
  assign n33951 = ~n26115 ;
  assign n26116 = x[59] & n33951 ;
  assign n26117 = n30638 & n26115 ;
  assign n26118 = n26116 | n26117 ;
  assign n26119 = n26111 | n26118 ;
  assign n26120 = n26111 & n26118 ;
  assign n33952 = ~n26120 ;
  assign n26121 = n26119 & n33952 ;
  assign n26122 = n25977 | n25987 ;
  assign n26123 = n26121 | n26122 ;
  assign n26124 = n26121 & n26122 ;
  assign n33953 = ~n26124 ;
  assign n26125 = n26123 & n33953 ;
  assign n26126 = n26090 | n26125 ;
  assign n26127 = n26090 & n26125 ;
  assign n33954 = ~n26127 ;
  assign n26128 = n26126 & n33954 ;
  assign n26129 = n26083 & n26128 ;
  assign n26130 = n26083 | n26128 ;
  assign n33955 = ~n26129 ;
  assign n26131 = n33955 & n26130 ;
  assign n1691 = n784 & n1690 ;
  assign n1555 = x[116] & n1551 ;
  assign n1628 = x[117] & n1616 ;
  assign n26132 = n1555 | n1628 ;
  assign n26133 = x[118] & n1547 ;
  assign n26134 = n26132 | n26133 ;
  assign n26135 = n1691 | n26134 ;
  assign n33956 = ~n26135 ;
  assign n26136 = x[53] & n33956 ;
  assign n26137 = n30125 & n26135 ;
  assign n26138 = n26136 | n26137 ;
  assign n33957 = ~n26138 ;
  assign n26139 = n26131 & n33957 ;
  assign n33958 = ~n26131 ;
  assign n26140 = n33958 & n26138 ;
  assign n26141 = n26139 | n26140 ;
  assign n26142 = n26080 | n26141 ;
  assign n26143 = n26080 & n26141 ;
  assign n33959 = ~n26143 ;
  assign n26144 = n26142 & n33959 ;
  assign n26145 = n26078 | n26144 ;
  assign n26146 = n26078 & n26144 ;
  assign n33960 = ~n26146 ;
  assign n26147 = n26145 & n33960 ;
  assign n26148 = n26071 | n26147 ;
  assign n26149 = n26071 & n26147 ;
  assign n33961 = ~n26149 ;
  assign n26150 = n26148 & n33961 ;
  assign n5842 = n2321 & n5838 ;
  assign n2221 = x[122] & n2179 ;
  assign n2264 = x[123] & n2244 ;
  assign n26151 = n2221 | n2264 ;
  assign n26152 = x[124] & n2175 ;
  assign n26153 = n26151 | n26152 ;
  assign n26154 = n5842 | n26153 ;
  assign n33962 = ~n26154 ;
  assign n26155 = x[47] & n33962 ;
  assign n26156 = n29621 & n26154 ;
  assign n26157 = n26155 | n26156 ;
  assign n26158 = n26150 | n26157 ;
  assign n26159 = n26150 & n26157 ;
  assign n33963 = ~n26159 ;
  assign n26160 = n26158 & n33963 ;
  assign n33964 = ~n26032 ;
  assign n26161 = n33964 & n26039 ;
  assign n26162 = n26031 | n26161 ;
  assign n33965 = ~n26162 ;
  assign n26163 = n26160 & n33965 ;
  assign n33966 = ~n26160 ;
  assign n26164 = n33966 & n26162 ;
  assign n26165 = n26163 | n26164 ;
  assign n5638 = n2635 & n5629 ;
  assign n2535 = x[125] & n2492 ;
  assign n2619 = x[126] & n2557 ;
  assign n26166 = n2535 | n2619 ;
  assign n26167 = x[127] & n2488 ;
  assign n26168 = n26166 | n26167 ;
  assign n26169 = n5638 | n26168 ;
  assign n33967 = ~n26169 ;
  assign n26170 = x[44] & n33967 ;
  assign n26171 = n29400 & n26169 ;
  assign n26172 = n26170 | n26171 ;
  assign n26173 = n26165 | n26172 ;
  assign n26174 = n26165 & n26172 ;
  assign n33968 = ~n26174 ;
  assign n26175 = n26173 & n33968 ;
  assign n33969 = ~n26048 ;
  assign n26176 = n33969 & n26055 ;
  assign n26177 = n26047 | n26176 ;
  assign n26178 = n26175 | n26177 ;
  assign n26179 = n26175 & n26177 ;
  assign n33970 = ~n26179 ;
  assign n26180 = n26178 & n33970 ;
  assign n33971 = ~n26058 ;
  assign n26059 = n25950 & n33971 ;
  assign n26181 = n25949 | n26059 ;
  assign n26182 = n26180 | n26181 ;
  assign n26183 = n26180 & n26181 ;
  assign n33972 = ~n26183 ;
  assign n26184 = n26182 & n33972 ;
  assign n26185 = n26069 & n26184 ;
  assign n26186 = n26069 | n26184 ;
  assign n33973 = ~n26185 ;
  assign n234 = n33973 & n26186 ;
  assign n33974 = ~n26150 ;
  assign n26188 = n33974 & n26157 ;
  assign n26189 = n26164 | n26188 ;
  assign n6195 = n2635 & n6186 ;
  assign n2552 = x[126] & n2492 ;
  assign n26190 = x[127] & n2557 ;
  assign n26191 = n2552 | n26190 ;
  assign n26192 = n6195 | n26191 ;
  assign n33975 = ~n26192 ;
  assign n26193 = x[44] & n33975 ;
  assign n26194 = n29400 & n26192 ;
  assign n26195 = n26193 | n26194 ;
  assign n26196 = n26189 | n26195 ;
  assign n26197 = n26189 & n26195 ;
  assign n33976 = ~n26197 ;
  assign n26198 = n26196 & n33976 ;
  assign n2344 = n642 & n2321 ;
  assign n2240 = x[123] & n2179 ;
  assign n2266 = x[124] & n2244 ;
  assign n26199 = n2240 | n2266 ;
  assign n26200 = x[125] & n2175 ;
  assign n26201 = n26199 | n26200 ;
  assign n26202 = n2344 | n26201 ;
  assign n26203 = x[47] | n26202 ;
  assign n26204 = x[47] & n26202 ;
  assign n33977 = ~n26204 ;
  assign n26205 = n26203 & n33977 ;
  assign n33978 = ~n26144 ;
  assign n26206 = n26078 & n33978 ;
  assign n33979 = ~n26147 ;
  assign n26207 = n26071 & n33979 ;
  assign n26208 = n26206 | n26207 ;
  assign n33980 = ~n26141 ;
  assign n26209 = n26080 & n33980 ;
  assign n26210 = n26140 | n26209 ;
  assign n33981 = ~n26096 ;
  assign n26211 = n33981 & n26103 ;
  assign n26212 = n26110 | n26211 ;
  assign n297 = x[106] & n27215 ;
  assign n832 = x[107] & n805 ;
  assign n26213 = n297 | n832 ;
  assign n26214 = n29184 & n25806 ;
  assign n26215 = n26095 | n26214 ;
  assign n26216 = n26213 | n26215 ;
  assign n26217 = n26213 & n26215 ;
  assign n33982 = ~n26217 ;
  assign n26218 = n26216 & n33982 ;
  assign n888 = x[110] & n881 ;
  assign n26219 = x[108] & n900 ;
  assign n26220 = x[109] & n949 ;
  assign n26221 = n26219 | n26220 ;
  assign n26222 = n888 | n26221 ;
  assign n26223 = n1006 & n3615 ;
  assign n26224 = n26222 | n26223 ;
  assign n26225 = n30886 & n26224 ;
  assign n33983 = ~n26224 ;
  assign n26226 = x[62] & n33983 ;
  assign n26227 = n26225 | n26226 ;
  assign n33984 = ~n26227 ;
  assign n26228 = n26218 & n33984 ;
  assign n33985 = ~n26218 ;
  assign n26229 = n33985 & n26227 ;
  assign n26230 = n26228 | n26229 ;
  assign n26231 = n26212 | n26230 ;
  assign n26232 = n26212 & n26230 ;
  assign n33986 = ~n26232 ;
  assign n26233 = n26231 & n33986 ;
  assign n4088 = n1217 & n4087 ;
  assign n1085 = x[111] & n1079 ;
  assign n1171 = x[112] & n1144 ;
  assign n26234 = n1085 | n1171 ;
  assign n26235 = x[113] & n1075 ;
  assign n26236 = n26234 | n26235 ;
  assign n26237 = n4088 | n26236 ;
  assign n33987 = ~n26237 ;
  assign n26238 = x[59] & n33987 ;
  assign n26239 = n30638 & n26237 ;
  assign n26240 = n26238 | n26239 ;
  assign n26241 = n26233 | n26240 ;
  assign n26242 = n26233 & n26240 ;
  assign n33988 = ~n26242 ;
  assign n26243 = n26241 & n33988 ;
  assign n33989 = ~n26111 ;
  assign n26244 = n33989 & n26118 ;
  assign n33990 = ~n26121 ;
  assign n26245 = n33990 & n26122 ;
  assign n26246 = n26244 | n26245 ;
  assign n33991 = ~n26246 ;
  assign n26247 = n26243 & n33991 ;
  assign n33992 = ~n26243 ;
  assign n26248 = n33992 & n26246 ;
  assign n26249 = n26247 | n26248 ;
  assign n4704 = n1457 & n4702 ;
  assign n1326 = x[114] & n1319 ;
  assign n1400 = x[115] & n1384 ;
  assign n26250 = n1326 | n1400 ;
  assign n26251 = x[116] & n1315 ;
  assign n26252 = n26250 | n26251 ;
  assign n26253 = n4704 | n26252 ;
  assign n33993 = ~n26253 ;
  assign n26254 = x[56] & n33993 ;
  assign n26255 = n30379 & n26253 ;
  assign n26256 = n26254 | n26255 ;
  assign n26257 = n26249 | n26256 ;
  assign n26258 = n26249 & n26256 ;
  assign n33994 = ~n26258 ;
  assign n26259 = n26257 & n33994 ;
  assign n33995 = ~n26125 ;
  assign n26260 = n26090 & n33995 ;
  assign n33996 = ~n26128 ;
  assign n26261 = n26083 & n33996 ;
  assign n26262 = n26260 | n26261 ;
  assign n33997 = ~n26262 ;
  assign n26263 = n26259 & n33997 ;
  assign n33998 = ~n26259 ;
  assign n26264 = n33998 & n26262 ;
  assign n26265 = n26263 | n26264 ;
  assign n5059 = n1690 & n5047 ;
  assign n1552 = x[117] & n1551 ;
  assign n1620 = x[118] & n1616 ;
  assign n26266 = n1552 | n1620 ;
  assign n26267 = x[119] & n1547 ;
  assign n26268 = n26266 | n26267 ;
  assign n26269 = n5059 | n26268 ;
  assign n33999 = ~n26269 ;
  assign n26270 = x[53] & n33999 ;
  assign n26271 = n30125 & n26269 ;
  assign n26272 = n26270 | n26271 ;
  assign n26273 = n26265 | n26272 ;
  assign n26274 = n26265 & n26272 ;
  assign n34000 = ~n26274 ;
  assign n26275 = n26273 & n34000 ;
  assign n26276 = n26210 & n26275 ;
  assign n26277 = n26210 | n26275 ;
  assign n34001 = ~n26276 ;
  assign n26278 = n34001 & n26277 ;
  assign n5028 = n2007 & n5022 ;
  assign n1882 = x[120] & n1866 ;
  assign n1933 = x[121] & n1931 ;
  assign n26279 = n1882 | n1933 ;
  assign n26280 = x[122] & n1862 ;
  assign n26281 = n26279 | n26280 ;
  assign n26282 = n5028 | n26281 ;
  assign n34002 = ~n26282 ;
  assign n26283 = x[50] & n34002 ;
  assign n26284 = n29865 & n26282 ;
  assign n26285 = n26283 | n26284 ;
  assign n26286 = n26278 | n26285 ;
  assign n26287 = n26278 & n26285 ;
  assign n34003 = ~n26287 ;
  assign n26288 = n26286 & n34003 ;
  assign n26289 = n26208 | n26288 ;
  assign n26290 = n26208 & n26288 ;
  assign n34004 = ~n26290 ;
  assign n26291 = n26289 & n34004 ;
  assign n26292 = n26205 & n26291 ;
  assign n26293 = n26205 | n26291 ;
  assign n34005 = ~n26292 ;
  assign n26294 = n34005 & n26293 ;
  assign n26295 = n26198 & n26294 ;
  assign n26296 = n26198 | n26294 ;
  assign n34006 = ~n26295 ;
  assign n26297 = n34006 & n26296 ;
  assign n34007 = ~n26165 ;
  assign n26298 = n34007 & n26172 ;
  assign n34008 = ~n26175 ;
  assign n26299 = n34008 & n26177 ;
  assign n26300 = n26298 | n26299 ;
  assign n34009 = ~n26300 ;
  assign n26301 = n26297 & n34009 ;
  assign n34010 = ~n26297 ;
  assign n26302 = n34010 & n26300 ;
  assign n26303 = n26301 | n26302 ;
  assign n34011 = ~n26180 ;
  assign n26304 = n34011 & n26181 ;
  assign n34012 = ~n26304 ;
  assign n26305 = n26186 & n34012 ;
  assign n26306 = n26303 | n26305 ;
  assign n26307 = n26303 & n26305 ;
  assign n34013 = ~n26307 ;
  assign n235 = n26306 & n34013 ;
  assign n34014 = ~n26302 ;
  assign n26309 = n34014 & n26306 ;
  assign n34015 = ~n26294 ;
  assign n26310 = n26198 & n34015 ;
  assign n26311 = n26197 | n26310 ;
  assign n34016 = ~n26288 ;
  assign n26312 = n26208 & n34016 ;
  assign n34017 = ~n26291 ;
  assign n26313 = n26205 & n34017 ;
  assign n26314 = n26312 | n26313 ;
  assign n2556 = x[127] & n2492 ;
  assign n5370 = n2635 & n5360 ;
  assign n26315 = n2556 | n5370 ;
  assign n34018 = ~n26315 ;
  assign n26316 = x[44] & n34018 ;
  assign n26317 = n29400 & n26315 ;
  assign n26318 = n26316 | n26317 ;
  assign n26319 = n26314 | n26318 ;
  assign n26320 = n26314 & n26318 ;
  assign n34019 = ~n26320 ;
  assign n26321 = n26319 & n34019 ;
  assign n34020 = ~n26265 ;
  assign n26322 = n34020 & n26272 ;
  assign n26323 = n26264 | n26322 ;
  assign n4689 = n1690 & n4678 ;
  assign n1587 = x[118] & n1551 ;
  assign n1649 = x[119] & n1616 ;
  assign n26376 = n1587 | n1649 ;
  assign n26377 = x[120] & n1547 ;
  assign n26378 = n26376 | n26377 ;
  assign n26379 = n4689 | n26378 ;
  assign n26380 = x[53] | n26379 ;
  assign n26381 = x[53] & n26379 ;
  assign n34021 = ~n26381 ;
  assign n26382 = n26380 & n34021 ;
  assign n34022 = ~n26249 ;
  assign n26324 = n34022 & n26256 ;
  assign n26325 = n26248 | n26324 ;
  assign n1458 = n797 & n1457 ;
  assign n1344 = x[115] & n1319 ;
  assign n1439 = x[116] & n1384 ;
  assign n26362 = n1344 | n1439 ;
  assign n26363 = x[117] & n1315 ;
  assign n26364 = n26362 | n26363 ;
  assign n26365 = n1458 | n26364 ;
  assign n26366 = x[56] | n26365 ;
  assign n26367 = x[56] & n26365 ;
  assign n34023 = ~n26367 ;
  assign n26368 = n26366 & n34023 ;
  assign n34024 = ~n26230 ;
  assign n26326 = n26212 & n34024 ;
  assign n34025 = ~n26233 ;
  assign n26327 = n34025 & n26240 ;
  assign n26328 = n26326 | n26327 ;
  assign n4281 = n1217 & n4276 ;
  assign n1084 = x[112] & n1079 ;
  assign n1152 = x[113] & n1144 ;
  assign n26349 = n1084 | n1152 ;
  assign n26350 = x[114] & n1075 ;
  assign n26351 = n26349 | n26350 ;
  assign n26352 = n4281 | n26351 ;
  assign n26353 = x[59] | n26352 ;
  assign n26354 = x[59] & n26352 ;
  assign n34026 = ~n26354 ;
  assign n26355 = n26353 & n34026 ;
  assign n34027 = ~n26213 ;
  assign n26329 = n34027 & n26215 ;
  assign n26330 = n26229 | n26329 ;
  assign n298 = x[107] & n27215 ;
  assign n817 = x[108] & n805 ;
  assign n26331 = n298 | n817 ;
  assign n26332 = n26213 | n26331 ;
  assign n26333 = n26213 & n26331 ;
  assign n34028 = ~n26333 ;
  assign n26334 = n26332 & n34028 ;
  assign n883 = x[111] & n881 ;
  assign n26335 = x[109] & n900 ;
  assign n26336 = x[110] & n949 ;
  assign n26337 = n26335 | n26336 ;
  assign n26338 = n883 | n26337 ;
  assign n26339 = n1006 & n4246 ;
  assign n26340 = n26338 | n26339 ;
  assign n26341 = n30886 & n26340 ;
  assign n34029 = ~n26340 ;
  assign n26342 = x[62] & n34029 ;
  assign n26343 = n26341 | n26342 ;
  assign n26344 = n26334 | n26343 ;
  assign n26345 = n26334 & n26343 ;
  assign n34030 = ~n26345 ;
  assign n26346 = n26344 & n34030 ;
  assign n26347 = n26330 | n26346 ;
  assign n26348 = n26330 & n26346 ;
  assign n34031 = ~n26348 ;
  assign n26356 = n26347 & n34031 ;
  assign n34032 = ~n26356 ;
  assign n26357 = n26355 & n34032 ;
  assign n34033 = ~n26355 ;
  assign n26358 = n26347 & n34033 ;
  assign n26359 = n34031 & n26358 ;
  assign n26360 = n26357 | n26359 ;
  assign n26361 = n26328 & n26360 ;
  assign n26369 = n26328 | n26360 ;
  assign n34034 = ~n26361 ;
  assign n26370 = n34034 & n26369 ;
  assign n34035 = ~n26370 ;
  assign n26371 = n26368 & n34035 ;
  assign n34036 = ~n26368 ;
  assign n26372 = n34036 & n26369 ;
  assign n26373 = n34034 & n26372 ;
  assign n26374 = n26371 | n26373 ;
  assign n26375 = n26325 & n26374 ;
  assign n26383 = n26325 | n26374 ;
  assign n34037 = ~n26375 ;
  assign n26384 = n34037 & n26383 ;
  assign n34038 = ~n26384 ;
  assign n26385 = n26382 & n34038 ;
  assign n34039 = ~n26382 ;
  assign n26386 = n34039 & n26383 ;
  assign n26387 = n34037 & n26386 ;
  assign n26388 = n26385 | n26387 ;
  assign n34040 = ~n26323 ;
  assign n26389 = n34040 & n26388 ;
  assign n34041 = ~n26388 ;
  assign n26390 = n26323 & n34041 ;
  assign n26391 = n26389 | n26390 ;
  assign n5430 = n2007 & n5417 ;
  assign n1867 = x[121] & n1866 ;
  assign n1932 = x[122] & n1931 ;
  assign n26392 = n1867 | n1932 ;
  assign n26393 = x[123] & n1862 ;
  assign n26394 = n26392 | n26393 ;
  assign n26395 = n5430 | n26394 ;
  assign n34042 = ~n26395 ;
  assign n26396 = x[50] & n34042 ;
  assign n26397 = n29865 & n26395 ;
  assign n26398 = n26396 | n26397 ;
  assign n26399 = n26391 | n26398 ;
  assign n26400 = n26391 & n26398 ;
  assign n34043 = ~n26400 ;
  assign n26401 = n26399 & n34043 ;
  assign n34044 = ~n26278 ;
  assign n26402 = n34044 & n26285 ;
  assign n34045 = ~n26275 ;
  assign n26403 = n26210 & n34045 ;
  assign n26404 = n26402 | n26403 ;
  assign n34046 = ~n26404 ;
  assign n26405 = n26401 & n34046 ;
  assign n34047 = ~n26401 ;
  assign n26406 = n34047 & n26404 ;
  assign n26407 = n26405 | n26406 ;
  assign n5389 = n2321 & n5388 ;
  assign n2226 = x[124] & n2179 ;
  assign n2304 = x[125] & n2244 ;
  assign n26408 = n2226 | n2304 ;
  assign n26409 = x[126] & n2175 ;
  assign n26410 = n26408 | n26409 ;
  assign n26411 = n5389 | n26410 ;
  assign n34048 = ~n26411 ;
  assign n26412 = x[47] & n34048 ;
  assign n26413 = n29621 & n26411 ;
  assign n26414 = n26412 | n26413 ;
  assign n34049 = ~n26414 ;
  assign n26415 = n26407 & n34049 ;
  assign n34050 = ~n26407 ;
  assign n26416 = n34050 & n26414 ;
  assign n26417 = n26415 | n26416 ;
  assign n26419 = n26321 & n26417 ;
  assign n26420 = n26321 | n26417 ;
  assign n34051 = ~n26419 ;
  assign n26421 = n34051 & n26420 ;
  assign n34052 = ~n26311 ;
  assign n26422 = n34052 & n26421 ;
  assign n34053 = ~n26421 ;
  assign n26423 = n26311 & n34053 ;
  assign n26424 = n26422 | n26423 ;
  assign n26425 = n26309 & n26424 ;
  assign n26426 = n26309 | n26424 ;
  assign n34054 = ~n26425 ;
  assign n236 = n34054 & n26426 ;
  assign n34055 = ~n26423 ;
  assign n26428 = n34055 & n26426 ;
  assign n34056 = ~n26391 ;
  assign n26429 = n34056 & n26398 ;
  assign n26430 = n26390 | n26429 ;
  assign n5847 = n2007 & n5838 ;
  assign n1913 = x[122] & n1866 ;
  assign n1991 = x[123] & n1931 ;
  assign n26431 = n1913 | n1991 ;
  assign n26432 = x[124] & n1862 ;
  assign n26433 = n26431 | n26432 ;
  assign n26434 = n5847 | n26433 ;
  assign n26435 = x[50] | n26434 ;
  assign n26436 = x[50] & n26434 ;
  assign n34057 = ~n26436 ;
  assign n26437 = n26435 & n34057 ;
  assign n34058 = ~n26374 ;
  assign n26438 = n26325 & n34058 ;
  assign n26439 = n26385 | n26438 ;
  assign n4997 = n1690 & n4985 ;
  assign n1554 = x[119] & n1551 ;
  assign n1619 = x[120] & n1616 ;
  assign n26440 = n1554 | n1619 ;
  assign n26441 = x[121] & n1547 ;
  assign n26442 = n26440 | n26441 ;
  assign n26443 = n4997 | n26442 ;
  assign n34059 = ~n26443 ;
  assign n26444 = x[53] & n34059 ;
  assign n26445 = n30125 & n26443 ;
  assign n26446 = n26444 | n26445 ;
  assign n34060 = ~n26360 ;
  assign n26447 = n26328 & n34060 ;
  assign n26448 = n26371 | n26447 ;
  assign n1461 = n784 & n1457 ;
  assign n1323 = x[116] & n1319 ;
  assign n1407 = x[117] & n1384 ;
  assign n26449 = n1323 | n1407 ;
  assign n26450 = x[118] & n1315 ;
  assign n26451 = n26449 | n26450 ;
  assign n26452 = n1461 | n26451 ;
  assign n26453 = x[56] | n26452 ;
  assign n26454 = x[56] & n26452 ;
  assign n34061 = ~n26454 ;
  assign n26455 = n26453 & n34061 ;
  assign n34062 = ~n26346 ;
  assign n26456 = n26330 & n34062 ;
  assign n26457 = n26357 | n26456 ;
  assign n26458 = n34027 & n26331 ;
  assign n34063 = ~n26334 ;
  assign n26459 = n34063 & n26343 ;
  assign n26460 = n26458 | n26459 ;
  assign n299 = x[108] & n27215 ;
  assign n816 = x[109] & n805 ;
  assign n26461 = n299 | n816 ;
  assign n34064 = ~n26461 ;
  assign n26462 = x[44] & n34064 ;
  assign n26463 = n29400 & n26461 ;
  assign n26464 = n26462 | n26463 ;
  assign n26465 = n26213 | n26464 ;
  assign n26467 = n26213 & n26464 ;
  assign n34065 = ~n26467 ;
  assign n26468 = n26465 & n34065 ;
  assign n34066 = ~n26460 ;
  assign n26469 = n34066 & n26468 ;
  assign n34067 = ~n26468 ;
  assign n26470 = n26460 & n34067 ;
  assign n26471 = n26469 | n26470 ;
  assign n4454 = n1006 & n4442 ;
  assign n904 = x[110] & n900 ;
  assign n991 = x[111] & n949 ;
  assign n26472 = n904 | n991 ;
  assign n26473 = x[112] & n881 ;
  assign n26474 = n26472 | n26473 ;
  assign n26475 = n4454 | n26474 ;
  assign n34068 = ~n26475 ;
  assign n26476 = x[62] & n34068 ;
  assign n26477 = n30886 & n26475 ;
  assign n26478 = n26476 | n26477 ;
  assign n34069 = ~n26478 ;
  assign n26479 = n26471 & n34069 ;
  assign n34070 = ~n26471 ;
  assign n26480 = n34070 & n26478 ;
  assign n26481 = n26479 | n26480 ;
  assign n4485 = n1217 & n4474 ;
  assign n1141 = x[113] & n1079 ;
  assign n1185 = x[114] & n1144 ;
  assign n26482 = n1141 | n1185 ;
  assign n26483 = x[115] & n1075 ;
  assign n26484 = n26482 | n26483 ;
  assign n26485 = n4485 | n26484 ;
  assign n34071 = ~n26485 ;
  assign n26486 = x[59] & n34071 ;
  assign n26487 = n30638 & n26485 ;
  assign n26488 = n26486 | n26487 ;
  assign n34072 = ~n26488 ;
  assign n26489 = n26481 & n34072 ;
  assign n34073 = ~n26481 ;
  assign n26490 = n34073 & n26488 ;
  assign n26491 = n26489 | n26490 ;
  assign n26492 = n26457 | n26491 ;
  assign n26494 = n26457 & n26491 ;
  assign n34074 = ~n26494 ;
  assign n26495 = n26492 & n34074 ;
  assign n34075 = ~n26495 ;
  assign n26496 = n26455 & n34075 ;
  assign n34076 = ~n26455 ;
  assign n26497 = n34076 & n26495 ;
  assign n26498 = n26496 | n26497 ;
  assign n26499 = n26448 | n26498 ;
  assign n26500 = n26448 & n26498 ;
  assign n34077 = ~n26500 ;
  assign n26501 = n26499 & n34077 ;
  assign n26502 = n26446 | n26501 ;
  assign n26503 = n26446 & n26501 ;
  assign n34078 = ~n26503 ;
  assign n26504 = n26502 & n34078 ;
  assign n26505 = n26439 | n26504 ;
  assign n26506 = n26439 & n26504 ;
  assign n34079 = ~n26506 ;
  assign n26507 = n26505 & n34079 ;
  assign n34080 = ~n26507 ;
  assign n26508 = n26437 & n34080 ;
  assign n34081 = ~n26437 ;
  assign n26509 = n34081 & n26507 ;
  assign n26510 = n26508 | n26509 ;
  assign n26511 = n26430 | n26510 ;
  assign n26512 = n26430 & n26510 ;
  assign n34082 = ~n26512 ;
  assign n26513 = n26511 & n34082 ;
  assign n5634 = n2321 & n5629 ;
  assign n2241 = x[125] & n2179 ;
  assign n2306 = x[126] & n2244 ;
  assign n26514 = n2241 | n2306 ;
  assign n26515 = x[127] & n2175 ;
  assign n26516 = n26514 | n26515 ;
  assign n26517 = n5634 | n26516 ;
  assign n34083 = ~n26517 ;
  assign n26518 = x[47] & n34083 ;
  assign n26519 = n29621 & n26517 ;
  assign n26520 = n26518 | n26519 ;
  assign n26521 = n26513 | n26520 ;
  assign n26522 = n26513 & n26520 ;
  assign n34084 = ~n26522 ;
  assign n26523 = n26521 & n34084 ;
  assign n26524 = n26406 | n26416 ;
  assign n26525 = n26523 | n26524 ;
  assign n26526 = n26523 & n26524 ;
  assign n34085 = ~n26526 ;
  assign n26527 = n26525 & n34085 ;
  assign n34086 = ~n26417 ;
  assign n26418 = n26321 & n34086 ;
  assign n26528 = n26320 | n26418 ;
  assign n26529 = n26527 | n26528 ;
  assign n26530 = n26527 & n26528 ;
  assign n34087 = ~n26530 ;
  assign n26531 = n26529 & n34087 ;
  assign n26532 = n26428 | n26531 ;
  assign n26533 = n26428 & n26531 ;
  assign n34088 = ~n26533 ;
  assign n237 = n26532 & n34088 ;
  assign n34089 = ~n26510 ;
  assign n26535 = n26430 & n34089 ;
  assign n26536 = n26508 | n26535 ;
  assign n6193 = n2321 & n6186 ;
  assign n2242 = x[126] & n2179 ;
  assign n26537 = x[127] & n2244 ;
  assign n26538 = n2242 | n26537 ;
  assign n26539 = n6193 | n26538 ;
  assign n34090 = ~n26539 ;
  assign n26540 = x[47] & n34090 ;
  assign n26541 = n29621 & n26539 ;
  assign n26542 = n26540 | n26541 ;
  assign n34091 = ~n26542 ;
  assign n26543 = n26536 & n34091 ;
  assign n34092 = ~n26536 ;
  assign n26544 = n34092 & n26542 ;
  assign n26545 = n26543 | n26544 ;
  assign n2026 = n642 & n2007 ;
  assign n1900 = x[123] & n1866 ;
  assign n1975 = x[124] & n1931 ;
  assign n26546 = n1900 | n1975 ;
  assign n26547 = x[125] & n1862 ;
  assign n26548 = n26546 | n26547 ;
  assign n26549 = n2026 | n26548 ;
  assign n26550 = x[50] | n26549 ;
  assign n26551 = x[50] & n26549 ;
  assign n34093 = ~n26551 ;
  assign n26552 = n26550 & n34093 ;
  assign n34094 = ~n26501 ;
  assign n26553 = n26446 & n34094 ;
  assign n34095 = ~n26504 ;
  assign n26554 = n26439 & n34095 ;
  assign n26555 = n26553 | n26554 ;
  assign n34096 = ~n26498 ;
  assign n26556 = n26448 & n34096 ;
  assign n26557 = n26496 | n26556 ;
  assign n34097 = ~n26491 ;
  assign n26493 = n26457 & n34097 ;
  assign n26558 = n26490 | n26493 ;
  assign n4713 = n1217 & n4702 ;
  assign n1102 = x[114] & n1079 ;
  assign n1162 = x[115] & n1144 ;
  assign n26577 = n1102 | n1162 ;
  assign n26578 = x[116] & n1075 ;
  assign n26579 = n26577 | n26578 ;
  assign n26580 = n4713 | n26579 ;
  assign n26581 = x[59] | n26580 ;
  assign n26582 = x[59] & n26580 ;
  assign n34098 = ~n26582 ;
  assign n26583 = n26581 & n34098 ;
  assign n26559 = n26470 | n26480 ;
  assign n300 = x[109] & n27215 ;
  assign n814 = x[110] & n805 ;
  assign n26560 = n300 | n814 ;
  assign n34099 = ~n26464 ;
  assign n26466 = n26213 & n34099 ;
  assign n26561 = n26463 | n26466 ;
  assign n26562 = n26560 | n26561 ;
  assign n26563 = n26560 & n26561 ;
  assign n34100 = ~n26563 ;
  assign n26564 = n26562 & n34100 ;
  assign n4097 = n1006 & n4087 ;
  assign n942 = x[111] & n900 ;
  assign n984 = x[112] & n949 ;
  assign n26565 = n942 | n984 ;
  assign n26566 = x[113] & n881 ;
  assign n26567 = n26565 | n26566 ;
  assign n26568 = n4097 | n26567 ;
  assign n34101 = ~n26568 ;
  assign n26569 = x[62] & n34101 ;
  assign n26570 = n30886 & n26568 ;
  assign n26571 = n26569 | n26570 ;
  assign n26572 = n26564 | n26571 ;
  assign n26573 = n26564 & n26571 ;
  assign n34102 = ~n26573 ;
  assign n26574 = n26572 & n34102 ;
  assign n26575 = n26559 | n26574 ;
  assign n26576 = n26559 & n26574 ;
  assign n34103 = ~n26576 ;
  assign n26584 = n26575 & n34103 ;
  assign n34104 = ~n26584 ;
  assign n26585 = n26583 & n34104 ;
  assign n34105 = ~n26583 ;
  assign n26586 = n26575 & n34105 ;
  assign n26587 = n34103 & n26586 ;
  assign n26588 = n26585 | n26587 ;
  assign n34106 = ~n26558 ;
  assign n26589 = n34106 & n26588 ;
  assign n34107 = ~n26588 ;
  assign n26590 = n26558 & n34107 ;
  assign n26591 = n26589 | n26590 ;
  assign n5060 = n1457 & n5047 ;
  assign n1320 = x[117] & n1319 ;
  assign n1388 = x[118] & n1384 ;
  assign n26592 = n1320 | n1388 ;
  assign n26593 = x[119] & n1315 ;
  assign n26594 = n26592 | n26593 ;
  assign n26595 = n5060 | n26594 ;
  assign n34108 = ~n26595 ;
  assign n26596 = x[56] & n34108 ;
  assign n26597 = n30379 & n26595 ;
  assign n26598 = n26596 | n26597 ;
  assign n26599 = n26591 | n26598 ;
  assign n26600 = n26591 & n26598 ;
  assign n34109 = ~n26600 ;
  assign n26601 = n26599 & n34109 ;
  assign n26602 = n26557 & n26601 ;
  assign n26603 = n26557 | n26601 ;
  assign n34110 = ~n26602 ;
  assign n26604 = n34110 & n26603 ;
  assign n5031 = n1690 & n5022 ;
  assign n1553 = x[120] & n1551 ;
  assign n1617 = x[121] & n1616 ;
  assign n26605 = n1553 | n1617 ;
  assign n26606 = x[122] & n1547 ;
  assign n26607 = n26605 | n26606 ;
  assign n26608 = n5031 | n26607 ;
  assign n34111 = ~n26608 ;
  assign n26609 = x[53] & n34111 ;
  assign n26610 = n30125 & n26608 ;
  assign n26611 = n26609 | n26610 ;
  assign n26612 = n26604 | n26611 ;
  assign n26613 = n26604 & n26611 ;
  assign n34112 = ~n26613 ;
  assign n26614 = n26612 & n34112 ;
  assign n26615 = n26555 | n26614 ;
  assign n26616 = n26555 & n26614 ;
  assign n34113 = ~n26616 ;
  assign n26617 = n26615 & n34113 ;
  assign n26618 = n26552 & n26617 ;
  assign n26619 = n26552 | n26617 ;
  assign n34114 = ~n26618 ;
  assign n26620 = n34114 & n26619 ;
  assign n26621 = n26545 & n26620 ;
  assign n26622 = n26545 | n26620 ;
  assign n34115 = ~n26621 ;
  assign n26623 = n34115 & n26622 ;
  assign n34116 = ~n26513 ;
  assign n26624 = n34116 & n26520 ;
  assign n34117 = ~n26523 ;
  assign n26625 = n34117 & n26524 ;
  assign n26626 = n26624 | n26625 ;
  assign n34118 = ~n26626 ;
  assign n26627 = n26623 & n34118 ;
  assign n34119 = ~n26623 ;
  assign n26628 = n34119 & n26626 ;
  assign n26629 = n26627 | n26628 ;
  assign n34120 = ~n26527 ;
  assign n26630 = n34120 & n26528 ;
  assign n34121 = ~n26630 ;
  assign n26631 = n26532 & n34121 ;
  assign n26632 = n26629 & n26631 ;
  assign n26633 = n26629 | n26631 ;
  assign n34122 = ~n26632 ;
  assign n238 = n34122 & n26633 ;
  assign n34123 = ~n26591 ;
  assign n26635 = n34123 & n26598 ;
  assign n26636 = n26590 | n26635 ;
  assign n4690 = n1457 & n4678 ;
  assign n1321 = x[118] & n1319 ;
  assign n1396 = x[119] & n1384 ;
  assign n26674 = n1321 | n1396 ;
  assign n26675 = x[120] & n1315 ;
  assign n26676 = n26674 | n26675 ;
  assign n26677 = n4690 | n26676 ;
  assign n26678 = x[56] | n26677 ;
  assign n26679 = x[56] & n26677 ;
  assign n34124 = ~n26679 ;
  assign n26680 = n26678 & n34124 ;
  assign n34125 = ~n26574 ;
  assign n26637 = n26559 & n34125 ;
  assign n26638 = n26585 | n26637 ;
  assign n1218 = n797 & n1217 ;
  assign n1083 = x[115] & n1079 ;
  assign n1151 = x[116] & n1144 ;
  assign n26639 = n1083 | n1151 ;
  assign n26640 = x[117] & n1075 ;
  assign n26641 = n26639 | n26640 ;
  assign n26642 = n1218 | n26641 ;
  assign n34126 = ~n26642 ;
  assign n26643 = x[59] & n34126 ;
  assign n26644 = n30638 & n26642 ;
  assign n26645 = n26643 | n26644 ;
  assign n34127 = ~n26560 ;
  assign n26649 = n34127 & n26561 ;
  assign n34128 = ~n26564 ;
  assign n26650 = n34128 & n26571 ;
  assign n26652 = n26649 | n26650 ;
  assign n301 = x[110] & n27215 ;
  assign n863 = x[111] & n805 ;
  assign n26646 = n301 | n863 ;
  assign n26648 = n34127 & n26646 ;
  assign n34129 = ~n26646 ;
  assign n26651 = n26560 & n34129 ;
  assign n26653 = n26648 | n26651 ;
  assign n26654 = n26652 & n26653 ;
  assign n34130 = ~n26648 ;
  assign n26655 = n34130 & n26652 ;
  assign n26656 = n26651 | n26655 ;
  assign n26657 = n26648 | n26656 ;
  assign n34131 = ~n26654 ;
  assign n26658 = n34131 & n26657 ;
  assign n4287 = n1006 & n4276 ;
  assign n938 = x[112] & n900 ;
  assign n992 = x[113] & n949 ;
  assign n26659 = n938 | n992 ;
  assign n26660 = x[114] & n881 ;
  assign n26661 = n26659 | n26660 ;
  assign n26662 = n4287 | n26661 ;
  assign n34132 = ~n26662 ;
  assign n26663 = x[62] & n34132 ;
  assign n26664 = n30886 & n26662 ;
  assign n26665 = n26663 | n26664 ;
  assign n26666 = n26658 | n26665 ;
  assign n26667 = n26658 & n26665 ;
  assign n34133 = ~n26667 ;
  assign n26668 = n26666 & n34133 ;
  assign n34134 = ~n26645 ;
  assign n26669 = n34134 & n26668 ;
  assign n34135 = ~n26668 ;
  assign n26670 = n26645 & n34135 ;
  assign n26671 = n26669 | n26670 ;
  assign n26672 = n26638 | n26671 ;
  assign n26673 = n26638 & n26671 ;
  assign n34136 = ~n26673 ;
  assign n26681 = n26672 & n34136 ;
  assign n34137 = ~n26681 ;
  assign n26682 = n26680 & n34137 ;
  assign n34138 = ~n26680 ;
  assign n26683 = n26672 & n34138 ;
  assign n26684 = n34136 & n26683 ;
  assign n26685 = n26682 | n26684 ;
  assign n34139 = ~n26636 ;
  assign n26686 = n34139 & n26685 ;
  assign n34140 = ~n26685 ;
  assign n26687 = n26636 & n34140 ;
  assign n26688 = n26686 | n26687 ;
  assign n5428 = n1690 & n5417 ;
  assign n1576 = x[121] & n1551 ;
  assign n1654 = x[122] & n1616 ;
  assign n26689 = n1576 | n1654 ;
  assign n26690 = x[123] & n1547 ;
  assign n26691 = n26689 | n26690 ;
  assign n26692 = n5428 | n26691 ;
  assign n34141 = ~n26692 ;
  assign n26693 = x[53] & n34141 ;
  assign n26694 = n30125 & n26692 ;
  assign n26695 = n26693 | n26694 ;
  assign n26696 = n26688 | n26695 ;
  assign n26697 = n26688 & n26695 ;
  assign n34142 = ~n26697 ;
  assign n26698 = n26696 & n34142 ;
  assign n34143 = ~n26604 ;
  assign n26699 = n34143 & n26611 ;
  assign n34144 = ~n26601 ;
  assign n26700 = n26557 & n34144 ;
  assign n26701 = n26699 | n26700 ;
  assign n34145 = ~n26701 ;
  assign n26702 = n26698 & n34145 ;
  assign n34146 = ~n26698 ;
  assign n26703 = n34146 & n26701 ;
  assign n26704 = n26702 | n26703 ;
  assign n5400 = n2007 & n5388 ;
  assign n1928 = x[124] & n1866 ;
  assign n1992 = x[125] & n1931 ;
  assign n26705 = n1928 | n1992 ;
  assign n26706 = x[126] & n1862 ;
  assign n26707 = n26705 | n26706 ;
  assign n26708 = n5400 | n26707 ;
  assign n34147 = ~n26708 ;
  assign n26709 = x[50] & n34147 ;
  assign n26710 = n29865 & n26708 ;
  assign n26711 = n26709 | n26710 ;
  assign n34148 = ~n26711 ;
  assign n26712 = n26704 & n34148 ;
  assign n34149 = ~n26704 ;
  assign n26713 = n34149 & n26711 ;
  assign n26714 = n26712 | n26713 ;
  assign n34150 = ~n26614 ;
  assign n26715 = n26555 & n34150 ;
  assign n34151 = ~n26617 ;
  assign n26716 = n26552 & n34151 ;
  assign n26717 = n26715 | n26716 ;
  assign n2243 = x[127] & n2179 ;
  assign n5368 = n2321 & n5360 ;
  assign n26718 = n2243 | n5368 ;
  assign n34152 = ~n26718 ;
  assign n26719 = x[47] & n34152 ;
  assign n26720 = n29621 & n26718 ;
  assign n26721 = n26719 | n26720 ;
  assign n26722 = n26717 | n26721 ;
  assign n26723 = n26717 & n26721 ;
  assign n34153 = ~n26723 ;
  assign n26724 = n26722 & n34153 ;
  assign n34154 = ~n26714 ;
  assign n26725 = n34154 & n26724 ;
  assign n34155 = ~n26724 ;
  assign n26726 = n26714 & n34155 ;
  assign n26727 = n26725 | n26726 ;
  assign n26728 = n26536 & n26542 ;
  assign n34156 = ~n26620 ;
  assign n26729 = n26545 & n34156 ;
  assign n26730 = n26728 | n26729 ;
  assign n34157 = ~n26730 ;
  assign n26731 = n26727 & n34157 ;
  assign n34158 = ~n26727 ;
  assign n26732 = n34158 & n26730 ;
  assign n26733 = n26731 | n26732 ;
  assign n34159 = ~n26628 ;
  assign n26734 = n34159 & n26633 ;
  assign n26735 = n26733 | n26734 ;
  assign n26736 = n26733 & n26734 ;
  assign n34160 = ~n26736 ;
  assign n239 = n26735 & n34160 ;
  assign n34161 = ~n26688 ;
  assign n26738 = n34161 & n26695 ;
  assign n26739 = n26687 | n26738 ;
  assign n5848 = n1690 & n5838 ;
  assign n1556 = x[122] & n1551 ;
  assign n1658 = x[123] & n1616 ;
  assign n26740 = n1556 | n1658 ;
  assign n26741 = x[124] & n1547 ;
  assign n26742 = n26740 | n26741 ;
  assign n26743 = n5848 | n26742 ;
  assign n26744 = x[53] | n26743 ;
  assign n26745 = x[53] & n26743 ;
  assign n34162 = ~n26745 ;
  assign n26746 = n26744 & n34162 ;
  assign n34163 = ~n26671 ;
  assign n26747 = n26638 & n34163 ;
  assign n26748 = n26682 | n26747 ;
  assign n4995 = n1457 & n4985 ;
  assign n1324 = x[119] & n1319 ;
  assign n1387 = x[120] & n1384 ;
  assign n26749 = n1324 | n1387 ;
  assign n26750 = x[121] & n1315 ;
  assign n26751 = n26749 | n26750 ;
  assign n26752 = n4995 | n26751 ;
  assign n34164 = ~n26752 ;
  assign n26753 = x[56] & n34164 ;
  assign n26754 = n30379 & n26752 ;
  assign n26755 = n26753 | n26754 ;
  assign n34165 = ~n26658 ;
  assign n26756 = n34165 & n26665 ;
  assign n26757 = n26670 | n26756 ;
  assign n4486 = n1006 & n4474 ;
  assign n931 = x[113] & n900 ;
  assign n993 = x[114] & n949 ;
  assign n26758 = n931 | n993 ;
  assign n26759 = x[115] & n881 ;
  assign n26760 = n26758 | n26759 ;
  assign n26761 = n4486 | n26760 ;
  assign n34166 = ~n26761 ;
  assign n26762 = x[62] & n34166 ;
  assign n26763 = n30886 & n26761 ;
  assign n26764 = n26762 | n26763 ;
  assign n302 = x[111] & n27215 ;
  assign n815 = x[112] & n805 ;
  assign n26765 = n302 | n815 ;
  assign n26647 = x[47] | n26646 ;
  assign n26766 = x[47] & n26646 ;
  assign n34167 = ~n26766 ;
  assign n26767 = n26647 & n34167 ;
  assign n34168 = ~n26765 ;
  assign n26768 = n34168 & n26767 ;
  assign n34169 = ~n26767 ;
  assign n26769 = n26765 & n34169 ;
  assign n26770 = n26768 | n26769 ;
  assign n26771 = n26764 | n26770 ;
  assign n26772 = n26764 & n26770 ;
  assign n34170 = ~n26772 ;
  assign n26773 = n26771 & n34170 ;
  assign n26774 = n26656 & n26773 ;
  assign n26775 = n26656 | n26773 ;
  assign n34171 = ~n26774 ;
  assign n26776 = n34171 & n26775 ;
  assign n1220 = n784 & n1217 ;
  assign n1139 = x[116] & n1079 ;
  assign n1150 = x[117] & n1144 ;
  assign n26777 = n1139 | n1150 ;
  assign n26778 = x[118] & n1075 ;
  assign n26779 = n26777 | n26778 ;
  assign n26780 = n1220 | n26779 ;
  assign n34172 = ~n26780 ;
  assign n26781 = x[59] & n34172 ;
  assign n26782 = n30638 & n26780 ;
  assign n26783 = n26781 | n26782 ;
  assign n34173 = ~n26783 ;
  assign n26784 = n26776 & n34173 ;
  assign n34174 = ~n26776 ;
  assign n26785 = n34174 & n26783 ;
  assign n26786 = n26784 | n26785 ;
  assign n26787 = n26757 | n26786 ;
  assign n26788 = n26757 & n26786 ;
  assign n34175 = ~n26788 ;
  assign n26789 = n26787 & n34175 ;
  assign n26790 = n26755 | n26789 ;
  assign n26791 = n26755 & n26789 ;
  assign n34176 = ~n26791 ;
  assign n26792 = n26790 & n34176 ;
  assign n26793 = n26748 | n26792 ;
  assign n26794 = n26748 & n26792 ;
  assign n34177 = ~n26794 ;
  assign n26795 = n26793 & n34177 ;
  assign n34178 = ~n26795 ;
  assign n26796 = n26746 & n34178 ;
  assign n34179 = ~n26746 ;
  assign n26797 = n34179 & n26795 ;
  assign n26798 = n26796 | n26797 ;
  assign n26799 = n26739 | n26798 ;
  assign n26800 = n26739 & n26798 ;
  assign n34180 = ~n26800 ;
  assign n26801 = n26799 & n34180 ;
  assign n5640 = n2007 & n5629 ;
  assign n1929 = x[125] & n1866 ;
  assign n1993 = x[126] & n1931 ;
  assign n26802 = n1929 | n1993 ;
  assign n26803 = x[127] & n1862 ;
  assign n26804 = n26802 | n26803 ;
  assign n26805 = n5640 | n26804 ;
  assign n34181 = ~n26805 ;
  assign n26806 = x[50] & n34181 ;
  assign n26807 = n29865 & n26805 ;
  assign n26808 = n26806 | n26807 ;
  assign n26809 = n26801 | n26808 ;
  assign n26810 = n26801 & n26808 ;
  assign n34182 = ~n26810 ;
  assign n26811 = n26809 & n34182 ;
  assign n26812 = n26703 | n26713 ;
  assign n26813 = n26811 | n26812 ;
  assign n26814 = n26811 & n26812 ;
  assign n34183 = ~n26814 ;
  assign n26815 = n26813 & n34183 ;
  assign n26816 = n26723 | n26725 ;
  assign n26817 = n26815 | n26816 ;
  assign n26818 = n26815 & n26816 ;
  assign n34184 = ~n26818 ;
  assign n26819 = n26817 & n34184 ;
  assign n34185 = ~n26732 ;
  assign n26820 = n34185 & n26735 ;
  assign n26821 = n26819 & n26820 ;
  assign n26822 = n26819 | n26820 ;
  assign n34186 = ~n26821 ;
  assign n240 = n34186 & n26822 ;
  assign n34187 = ~n26798 ;
  assign n26824 = n26739 & n34187 ;
  assign n26825 = n26796 | n26824 ;
  assign n1704 = n642 & n1690 ;
  assign n1582 = x[123] & n1551 ;
  assign n1676 = x[124] & n1616 ;
  assign n26826 = n1582 | n1676 ;
  assign n26827 = x[125] & n1547 ;
  assign n26828 = n26826 | n26827 ;
  assign n26829 = n1704 | n26828 ;
  assign n34188 = ~n26829 ;
  assign n26830 = x[53] & n34188 ;
  assign n26831 = n30125 & n26829 ;
  assign n26832 = n26830 | n26831 ;
  assign n34189 = ~n26789 ;
  assign n26833 = n26755 & n34189 ;
  assign n34190 = ~n26792 ;
  assign n26834 = n26748 & n34190 ;
  assign n26835 = n26833 | n26834 ;
  assign n5029 = n1457 & n5022 ;
  assign n1380 = x[120] & n1319 ;
  assign n1429 = x[121] & n1384 ;
  assign n26836 = n1380 | n1429 ;
  assign n26837 = x[122] & n1315 ;
  assign n26838 = n26836 | n26837 ;
  assign n26839 = n5029 | n26838 ;
  assign n26840 = x[56] | n26839 ;
  assign n26841 = x[56] & n26839 ;
  assign n34191 = ~n26841 ;
  assign n26842 = n26840 & n34191 ;
  assign n34192 = ~n26786 ;
  assign n26843 = n26757 & n34192 ;
  assign n26844 = n26785 | n26843 ;
  assign n5052 = n1217 & n5047 ;
  assign n1080 = x[117] & n1079 ;
  assign n1148 = x[118] & n1144 ;
  assign n26868 = n1080 | n1148 ;
  assign n26869 = x[119] & n1075 ;
  assign n26870 = n26868 | n26869 ;
  assign n26871 = n5052 | n26870 ;
  assign n26872 = x[59] | n26871 ;
  assign n26873 = x[59] & n26871 ;
  assign n34193 = ~n26873 ;
  assign n26874 = n26872 & n34193 ;
  assign n34194 = ~n26770 ;
  assign n26845 = n26764 & n34194 ;
  assign n34195 = ~n26773 ;
  assign n26846 = n26656 & n34195 ;
  assign n26847 = n26845 | n26846 ;
  assign n303 = x[112] & n27215 ;
  assign n856 = x[113] & n805 ;
  assign n26848 = n303 | n856 ;
  assign n26849 = n29621 & n26646 ;
  assign n26850 = n26769 | n26849 ;
  assign n34196 = ~n26850 ;
  assign n26851 = n26848 & n34196 ;
  assign n34197 = ~n26848 ;
  assign n26852 = n34197 & n26850 ;
  assign n26853 = n26851 | n26852 ;
  assign n894 = x[116] & n881 ;
  assign n26854 = x[114] & n900 ;
  assign n26855 = x[115] & n949 ;
  assign n26856 = n26854 | n26855 ;
  assign n26857 = n894 | n26856 ;
  assign n26858 = n1006 & n4702 ;
  assign n26859 = n26857 | n26858 ;
  assign n26860 = n30886 & n26859 ;
  assign n34198 = ~n26859 ;
  assign n26861 = x[62] & n34198 ;
  assign n26862 = n26860 | n26861 ;
  assign n26863 = n26853 | n26862 ;
  assign n26864 = n26853 & n26862 ;
  assign n34199 = ~n26864 ;
  assign n26865 = n26863 & n34199 ;
  assign n26866 = n26847 | n26865 ;
  assign n26867 = n26847 & n26865 ;
  assign n34200 = ~n26867 ;
  assign n26875 = n26866 & n34200 ;
  assign n34201 = ~n26875 ;
  assign n26876 = n26874 & n34201 ;
  assign n34202 = ~n26874 ;
  assign n26877 = n26866 & n34202 ;
  assign n26878 = n34200 & n26877 ;
  assign n26879 = n26876 | n26878 ;
  assign n26880 = n26844 & n26879 ;
  assign n26881 = n26844 | n26879 ;
  assign n34203 = ~n26880 ;
  assign n26882 = n34203 & n26881 ;
  assign n34204 = ~n26882 ;
  assign n26883 = n26842 & n34204 ;
  assign n34205 = ~n26842 ;
  assign n26884 = n34205 & n26882 ;
  assign n26885 = n26883 | n26884 ;
  assign n26886 = n26835 | n26885 ;
  assign n26887 = n26835 & n26885 ;
  assign n34206 = ~n26887 ;
  assign n26888 = n26886 & n34206 ;
  assign n34207 = ~n26888 ;
  assign n26889 = n26832 & n34207 ;
  assign n34208 = ~n26832 ;
  assign n26890 = n34208 & n26886 ;
  assign n26891 = n34206 & n26890 ;
  assign n26892 = n26889 | n26891 ;
  assign n34209 = ~n26892 ;
  assign n26893 = n26825 & n34209 ;
  assign n34210 = ~n26825 ;
  assign n26894 = n34210 & n26892 ;
  assign n26895 = n26893 | n26894 ;
  assign n6189 = n2007 & n6186 ;
  assign n1889 = x[126] & n1866 ;
  assign n26896 = x[127] & n1931 ;
  assign n26897 = n1889 | n26896 ;
  assign n26898 = n6189 | n26897 ;
  assign n34211 = ~n26898 ;
  assign n26899 = x[50] & n34211 ;
  assign n26900 = n29865 & n26898 ;
  assign n26901 = n26899 | n26900 ;
  assign n26902 = n26895 | n26901 ;
  assign n26903 = n26895 & n26901 ;
  assign n34212 = ~n26903 ;
  assign n26904 = n26902 & n34212 ;
  assign n34213 = ~n26801 ;
  assign n26905 = n34213 & n26808 ;
  assign n34214 = ~n26811 ;
  assign n26906 = n34214 & n26812 ;
  assign n26907 = n26905 | n26906 ;
  assign n34215 = ~n26907 ;
  assign n26908 = n26904 & n34215 ;
  assign n34216 = ~n26904 ;
  assign n26909 = n34216 & n26907 ;
  assign n26910 = n26908 | n26909 ;
  assign n34217 = ~n26815 ;
  assign n26911 = n34217 & n26816 ;
  assign n34218 = ~n26911 ;
  assign n26912 = n26822 & n34218 ;
  assign n26913 = n26910 | n26912 ;
  assign n26914 = n26910 & n26912 ;
  assign n34219 = ~n26914 ;
  assign n241 = n26913 & n34219 ;
  assign n34220 = ~n26865 ;
  assign n26916 = n26847 & n34220 ;
  assign n26917 = n26876 | n26916 ;
  assign n1009 = n797 & n1006 ;
  assign n943 = x[115] & n900 ;
  assign n987 = x[116] & n949 ;
  assign n26918 = n943 | n987 ;
  assign n26919 = x[117] & n881 ;
  assign n26920 = n26918 | n26919 ;
  assign n26921 = n1009 | n26920 ;
  assign n34221 = ~n26921 ;
  assign n26922 = x[62] & n34221 ;
  assign n26923 = n30886 & n26921 ;
  assign n26924 = n26922 | n26923 ;
  assign n304 = x[113] & n27215 ;
  assign n813 = x[114] & n805 ;
  assign n26925 = n304 | n813 ;
  assign n26926 = n26848 | n26925 ;
  assign n26927 = n26848 & n26925 ;
  assign n34222 = ~n26927 ;
  assign n26928 = n26926 & n34222 ;
  assign n34223 = ~n26924 ;
  assign n26929 = n34223 & n26928 ;
  assign n34224 = ~n26928 ;
  assign n26930 = n26924 & n34224 ;
  assign n26931 = n26929 | n26930 ;
  assign n34225 = ~n26853 ;
  assign n26932 = n34225 & n26862 ;
  assign n26933 = n26852 | n26932 ;
  assign n34226 = ~n26933 ;
  assign n26934 = n26931 & n34226 ;
  assign n34227 = ~n26931 ;
  assign n26935 = n34227 & n26933 ;
  assign n26936 = n26934 | n26935 ;
  assign n4683 = n1217 & n4678 ;
  assign n1100 = x[118] & n1079 ;
  assign n1145 = x[119] & n1144 ;
  assign n26937 = n1100 | n1145 ;
  assign n26938 = x[120] & n1075 ;
  assign n26939 = n26937 | n26938 ;
  assign n26940 = n4683 | n26939 ;
  assign n34228 = ~n26940 ;
  assign n26941 = x[59] & n34228 ;
  assign n26942 = n30638 & n26940 ;
  assign n26943 = n26941 | n26942 ;
  assign n26944 = n26936 | n26943 ;
  assign n26945 = n26936 & n26943 ;
  assign n34229 = ~n26945 ;
  assign n26946 = n26944 & n34229 ;
  assign n26947 = n26917 | n26946 ;
  assign n26948 = n26917 & n26946 ;
  assign n34230 = ~n26948 ;
  assign n26949 = n26947 & n34230 ;
  assign n5420 = n1457 & n5417 ;
  assign n1351 = x[121] & n1319 ;
  assign n1385 = x[122] & n1384 ;
  assign n26950 = n1351 | n1385 ;
  assign n26951 = x[123] & n1315 ;
  assign n26952 = n26950 | n26951 ;
  assign n26953 = n5420 | n26952 ;
  assign n34231 = ~n26953 ;
  assign n26954 = x[56] & n34231 ;
  assign n26955 = n30379 & n26953 ;
  assign n26956 = n26954 | n26955 ;
  assign n26957 = n26949 | n26956 ;
  assign n26958 = n26949 & n26956 ;
  assign n34232 = ~n26958 ;
  assign n26959 = n26957 & n34232 ;
  assign n34233 = ~n26879 ;
  assign n26960 = n26844 & n34233 ;
  assign n26961 = n26883 | n26960 ;
  assign n34234 = ~n26961 ;
  assign n26962 = n26959 & n34234 ;
  assign n34235 = ~n26959 ;
  assign n26963 = n34235 & n26961 ;
  assign n26964 = n26962 | n26963 ;
  assign n5401 = n1690 & n5388 ;
  assign n1613 = x[124] & n1551 ;
  assign n1677 = x[125] & n1616 ;
  assign n26965 = n1613 | n1677 ;
  assign n26966 = x[126] & n1547 ;
  assign n26967 = n26965 | n26966 ;
  assign n26968 = n5401 | n26967 ;
  assign n34236 = ~n26968 ;
  assign n26969 = x[53] & n34236 ;
  assign n26970 = n30125 & n26968 ;
  assign n26971 = n26969 | n26970 ;
  assign n26972 = n26964 | n26971 ;
  assign n26973 = n26964 & n26971 ;
  assign n34237 = ~n26973 ;
  assign n26974 = n26972 & n34237 ;
  assign n34238 = ~n26885 ;
  assign n26975 = n26835 & n34238 ;
  assign n26976 = n26889 | n26975 ;
  assign n1930 = x[127] & n1866 ;
  assign n5371 = n2007 & n5360 ;
  assign n26977 = n1930 | n5371 ;
  assign n34239 = ~n26977 ;
  assign n26978 = x[50] & n34239 ;
  assign n26979 = n29865 & n26977 ;
  assign n26980 = n26978 | n26979 ;
  assign n26981 = n26976 | n26980 ;
  assign n26982 = n26976 & n26980 ;
  assign n34240 = ~n26982 ;
  assign n26983 = n26981 & n34240 ;
  assign n34241 = ~n26974 ;
  assign n26984 = n34241 & n26983 ;
  assign n34242 = ~n26983 ;
  assign n26985 = n26974 & n34242 ;
  assign n26986 = n26984 | n26985 ;
  assign n34243 = ~n26895 ;
  assign n26987 = n34243 & n26901 ;
  assign n26988 = n26893 | n26987 ;
  assign n34244 = ~n26988 ;
  assign n26989 = n26986 & n34244 ;
  assign n34245 = ~n26986 ;
  assign n26990 = n34245 & n26988 ;
  assign n26991 = n26989 | n26990 ;
  assign n34246 = ~n26909 ;
  assign n26992 = n34246 & n26913 ;
  assign n26993 = n26991 & n26992 ;
  assign n26994 = n26991 | n26992 ;
  assign n34247 = ~n26993 ;
  assign n242 = n34247 & n26994 ;
  assign n34248 = ~n26946 ;
  assign n26996 = n26917 & n34248 ;
  assign n34249 = ~n26949 ;
  assign n26997 = n34249 & n26956 ;
  assign n26998 = n26996 | n26997 ;
  assign n5850 = n1457 & n5838 ;
  assign n1346 = x[122] & n1319 ;
  assign n1437 = x[123] & n1384 ;
  assign n26999 = n1346 | n1437 ;
  assign n27000 = x[124] & n1315 ;
  assign n27001 = n26999 | n27000 ;
  assign n27002 = n5850 | n27001 ;
  assign n27003 = x[56] | n27002 ;
  assign n27004 = x[56] & n27002 ;
  assign n34250 = ~n27004 ;
  assign n27005 = n27003 & n34250 ;
  assign n34251 = ~n26936 ;
  assign n27006 = n34251 & n26943 ;
  assign n27007 = n26935 | n27006 ;
  assign n4990 = n1217 & n4985 ;
  assign n1106 = x[119] & n1079 ;
  assign n1174 = x[120] & n1144 ;
  assign n27008 = n1106 | n1174 ;
  assign n27009 = x[121] & n1075 ;
  assign n27010 = n27008 | n27009 ;
  assign n27011 = n4990 | n27010 ;
  assign n34252 = ~n27011 ;
  assign n27012 = x[59] & n34252 ;
  assign n27013 = n30638 & n27011 ;
  assign n27014 = n27012 | n27013 ;
  assign n1007 = n784 & n1006 ;
  assign n926 = x[116] & n900 ;
  assign n994 = x[117] & n949 ;
  assign n27026 = n926 | n994 ;
  assign n27027 = x[118] & n881 ;
  assign n27028 = n27026 | n27027 ;
  assign n27029 = n1007 | n27028 ;
  assign n34253 = ~n27029 ;
  assign n27030 = x[62] & n34253 ;
  assign n27031 = n30886 & n27029 ;
  assign n27032 = n27030 | n27031 ;
  assign n27015 = n34197 & n26925 ;
  assign n27016 = n26930 | n27015 ;
  assign n305 = x[114] & n27215 ;
  assign n834 = x[115] & n805 ;
  assign n27017 = n305 | n834 ;
  assign n34254 = ~n27017 ;
  assign n27018 = x[50] & n34254 ;
  assign n27019 = n29865 & n27017 ;
  assign n27020 = n27018 | n27019 ;
  assign n34255 = ~n27020 ;
  assign n27021 = n26848 & n34255 ;
  assign n27022 = n34197 & n27020 ;
  assign n27023 = n27021 | n27022 ;
  assign n27024 = n27016 | n27023 ;
  assign n27025 = n27016 & n27023 ;
  assign n34256 = ~n27025 ;
  assign n27033 = n27024 & n34256 ;
  assign n34257 = ~n27033 ;
  assign n27034 = n27032 & n34257 ;
  assign n34258 = ~n27032 ;
  assign n27035 = n27024 & n34258 ;
  assign n27036 = n34256 & n27035 ;
  assign n27037 = n27034 | n27036 ;
  assign n27039 = n27014 & n27037 ;
  assign n27040 = n27014 | n27037 ;
  assign n34259 = ~n27039 ;
  assign n27041 = n34259 & n27040 ;
  assign n34260 = ~n27041 ;
  assign n27042 = n27007 & n34260 ;
  assign n34261 = ~n27007 ;
  assign n27043 = n34261 & n27040 ;
  assign n27044 = n34259 & n27043 ;
  assign n27045 = n27042 | n27044 ;
  assign n34262 = ~n27045 ;
  assign n27046 = n27005 & n34262 ;
  assign n34263 = ~n27005 ;
  assign n27047 = n34263 & n27045 ;
  assign n27048 = n27046 | n27047 ;
  assign n27049 = n26998 | n27048 ;
  assign n27050 = n26998 & n27048 ;
  assign n34264 = ~n27050 ;
  assign n27051 = n27049 & n34264 ;
  assign n5643 = n1690 & n5629 ;
  assign n1614 = x[125] & n1551 ;
  assign n1678 = x[126] & n1616 ;
  assign n27052 = n1614 | n1678 ;
  assign n27053 = x[127] & n1547 ;
  assign n27054 = n27052 | n27053 ;
  assign n27055 = n5643 | n27054 ;
  assign n34265 = ~n27055 ;
  assign n27056 = x[53] & n34265 ;
  assign n27057 = n30125 & n27055 ;
  assign n27058 = n27056 | n27057 ;
  assign n27059 = n27051 | n27058 ;
  assign n27060 = n27051 & n27058 ;
  assign n34266 = ~n27060 ;
  assign n27061 = n27059 & n34266 ;
  assign n34267 = ~n26964 ;
  assign n27062 = n34267 & n26971 ;
  assign n27063 = n26963 | n27062 ;
  assign n27064 = n27061 | n27063 ;
  assign n27065 = n27061 & n27063 ;
  assign n34268 = ~n27065 ;
  assign n27066 = n27064 & n34268 ;
  assign n27067 = n26982 | n26984 ;
  assign n27068 = n27066 | n27067 ;
  assign n27069 = n27066 & n27067 ;
  assign n34269 = ~n27069 ;
  assign n27070 = n27068 & n34269 ;
  assign n34270 = ~n26990 ;
  assign n27071 = n34270 & n26994 ;
  assign n27072 = n27070 | n27071 ;
  assign n27073 = n27070 & n27071 ;
  assign n34271 = ~n27073 ;
  assign n243 = n27072 & n34271 ;
  assign n34272 = ~n27048 ;
  assign n27075 = n26998 & n34272 ;
  assign n27076 = n27046 | n27075 ;
  assign n1468 = n642 & n1457 ;
  assign n1342 = x[123] & n1319 ;
  assign n1445 = x[124] & n1384 ;
  assign n27077 = n1342 | n1445 ;
  assign n27078 = x[125] & n1315 ;
  assign n27079 = n27077 | n27078 ;
  assign n27080 = n1468 | n27079 ;
  assign n34273 = ~n27080 ;
  assign n27081 = x[56] & n34273 ;
  assign n27082 = n30379 & n27080 ;
  assign n27083 = n27081 | n27082 ;
  assign n34274 = ~n27037 ;
  assign n27038 = n27014 & n34274 ;
  assign n27084 = n27038 | n27042 ;
  assign n5024 = n1217 & n5022 ;
  assign n1136 = x[120] & n1079 ;
  assign n1146 = x[121] & n1144 ;
  assign n27085 = n1136 | n1146 ;
  assign n27086 = x[122] & n1075 ;
  assign n27087 = n27085 | n27086 ;
  assign n27088 = n5024 | n27087 ;
  assign n34275 = ~n27088 ;
  assign n27089 = x[59] & n34275 ;
  assign n27090 = n30638 & n27088 ;
  assign n27091 = n27089 | n27090 ;
  assign n34276 = ~n27023 ;
  assign n27092 = n27016 & n34276 ;
  assign n27093 = n27034 | n27092 ;
  assign n306 = x[115] & n27215 ;
  assign n826 = x[116] & n805 ;
  assign n27094 = n306 | n826 ;
  assign n27095 = n27019 | n27021 ;
  assign n27096 = n27094 | n27095 ;
  assign n27097 = n27094 & n27095 ;
  assign n34277 = ~n27097 ;
  assign n27098 = n27096 & n34277 ;
  assign n5053 = n1006 & n5047 ;
  assign n945 = x[117] & n900 ;
  assign n974 = x[118] & n949 ;
  assign n27099 = n945 | n974 ;
  assign n27100 = x[119] & n881 ;
  assign n27101 = n27099 | n27100 ;
  assign n27102 = n5053 | n27101 ;
  assign n34278 = ~n27102 ;
  assign n27103 = x[62] & n34278 ;
  assign n27104 = n30886 & n27102 ;
  assign n27105 = n27103 | n27104 ;
  assign n27106 = n27098 | n27105 ;
  assign n27107 = n27098 & n27105 ;
  assign n34279 = ~n27107 ;
  assign n27108 = n27106 & n34279 ;
  assign n27109 = n27093 | n27108 ;
  assign n27110 = n27093 & n27108 ;
  assign n34280 = ~n27110 ;
  assign n27111 = n27109 & n34280 ;
  assign n27112 = n27091 | n27111 ;
  assign n27114 = n27091 & n27111 ;
  assign n34281 = ~n27114 ;
  assign n27115 = n27112 & n34281 ;
  assign n27116 = n27084 | n27115 ;
  assign n27117 = n27084 & n27115 ;
  assign n34282 = ~n27117 ;
  assign n27118 = n27116 & n34282 ;
  assign n34283 = ~n27118 ;
  assign n27119 = n27083 & n34283 ;
  assign n34284 = ~n27083 ;
  assign n27120 = n34284 & n27116 ;
  assign n27121 = n34282 & n27120 ;
  assign n27122 = n27119 | n27121 ;
  assign n34285 = ~n27122 ;
  assign n27123 = n27076 & n34285 ;
  assign n34286 = ~n27076 ;
  assign n27124 = n34286 & n27122 ;
  assign n27125 = n27123 | n27124 ;
  assign n6197 = n1690 & n6186 ;
  assign n1615 = x[126] & n1551 ;
  assign n27126 = x[127] & n1616 ;
  assign n27127 = n1615 | n27126 ;
  assign n27128 = n6197 | n27127 ;
  assign n34287 = ~n27128 ;
  assign n27129 = x[53] & n34287 ;
  assign n27130 = n30125 & n27128 ;
  assign n27131 = n27129 | n27130 ;
  assign n27132 = n27125 | n27131 ;
  assign n27133 = n27125 & n27131 ;
  assign n34288 = ~n27133 ;
  assign n27134 = n27132 & n34288 ;
  assign n34289 = ~n27051 ;
  assign n27135 = n34289 & n27058 ;
  assign n34290 = ~n27061 ;
  assign n27136 = n34290 & n27063 ;
  assign n27137 = n27135 | n27136 ;
  assign n34291 = ~n27137 ;
  assign n27138 = n27134 & n34291 ;
  assign n34292 = ~n27134 ;
  assign n27139 = n34292 & n27137 ;
  assign n27140 = n27138 | n27139 ;
  assign n34293 = ~n27066 ;
  assign n27141 = n34293 & n27067 ;
  assign n34294 = ~n27141 ;
  assign n27142 = n27072 & n34294 ;
  assign n27143 = n27140 & n27142 ;
  assign n27144 = n27140 | n27142 ;
  assign n34295 = ~n27143 ;
  assign n244 = n34295 & n27144 ;
  assign n34296 = ~n27111 ;
  assign n27113 = n27091 & n34296 ;
  assign n34297 = ~n27108 ;
  assign n27146 = n27093 & n34297 ;
  assign n27147 = n27113 | n27146 ;
  assign n34298 = ~n27094 ;
  assign n27148 = n34298 & n27095 ;
  assign n34299 = ~n27098 ;
  assign n27149 = n34299 & n27105 ;
  assign n27150 = n27148 | n27149 ;
  assign n307 = x[116] & n27215 ;
  assign n811 = x[117] & n805 ;
  assign n27151 = n307 | n811 ;
  assign n27153 = n34298 & n27151 ;
  assign n34300 = ~n27151 ;
  assign n27154 = n27094 & n34300 ;
  assign n27155 = n27153 | n27154 ;
  assign n27156 = n27150 & n27155 ;
  assign n34301 = ~n27153 ;
  assign n27157 = n27150 & n34301 ;
  assign n27158 = n27154 | n27157 ;
  assign n27159 = n27153 | n27158 ;
  assign n34302 = ~n27156 ;
  assign n27160 = n34302 & n27159 ;
  assign n4691 = n1006 & n4678 ;
  assign n946 = x[118] & n900 ;
  assign n995 = x[119] & n949 ;
  assign n27161 = n946 | n995 ;
  assign n27162 = x[120] & n881 ;
  assign n27163 = n27161 | n27162 ;
  assign n27164 = n4691 | n27163 ;
  assign n34303 = ~n27164 ;
  assign n27165 = x[62] & n34303 ;
  assign n27166 = n30886 & n27164 ;
  assign n27167 = n27165 | n27166 ;
  assign n34304 = ~n27167 ;
  assign n27168 = n27160 & n34304 ;
  assign n34305 = ~n27160 ;
  assign n27169 = n34305 & n27167 ;
  assign n27170 = n27168 | n27169 ;
  assign n5431 = n1217 & n5417 ;
  assign n1131 = x[121] & n1079 ;
  assign n1189 = x[122] & n1144 ;
  assign n27171 = n1131 | n1189 ;
  assign n27172 = x[123] & n1075 ;
  assign n27173 = n27171 | n27172 ;
  assign n27174 = n5431 | n27173 ;
  assign n34306 = ~n27174 ;
  assign n27175 = x[59] & n34306 ;
  assign n27176 = n30638 & n27174 ;
  assign n27177 = n27175 | n27176 ;
  assign n34307 = ~n27177 ;
  assign n27178 = n27170 & n34307 ;
  assign n34308 = ~n27170 ;
  assign n27179 = n34308 & n27177 ;
  assign n27180 = n27178 | n27179 ;
  assign n27181 = n27147 | n27180 ;
  assign n27182 = n27147 & n27180 ;
  assign n34309 = ~n27182 ;
  assign n27183 = n27181 & n34309 ;
  assign n5391 = n1457 & n5388 ;
  assign n1382 = x[124] & n1319 ;
  assign n1438 = x[125] & n1384 ;
  assign n27184 = n1382 | n1438 ;
  assign n27185 = x[126] & n1315 ;
  assign n27186 = n27184 | n27185 ;
  assign n27187 = n5391 | n27186 ;
  assign n34310 = ~n27187 ;
  assign n27188 = x[56] & n34310 ;
  assign n27189 = n30379 & n27187 ;
  assign n27190 = n27188 | n27189 ;
  assign n27191 = n27183 | n27190 ;
  assign n27192 = n27183 & n27190 ;
  assign n34311 = ~n27192 ;
  assign n27193 = n27191 & n34311 ;
  assign n34312 = ~n27115 ;
  assign n27194 = n27084 & n34312 ;
  assign n27195 = n27119 | n27194 ;
  assign n1592 = x[127] & n1551 ;
  assign n5372 = n1690 & n5360 ;
  assign n27196 = n1592 | n5372 ;
  assign n34313 = ~n27196 ;
  assign n27197 = x[53] & n34313 ;
  assign n27198 = n30125 & n27196 ;
  assign n27199 = n27197 | n27198 ;
  assign n27200 = n27195 | n27199 ;
  assign n27201 = n27195 & n27199 ;
  assign n34314 = ~n27201 ;
  assign n27202 = n27200 & n34314 ;
  assign n27203 = n27193 & n27202 ;
  assign n27205 = n27193 | n27202 ;
  assign n34315 = ~n27203 ;
  assign n27206 = n34315 & n27205 ;
  assign n34316 = ~n27125 ;
  assign n27207 = n34316 & n27131 ;
  assign n27208 = n27123 | n27207 ;
  assign n34317 = ~n27208 ;
  assign n27209 = n27206 & n34317 ;
  assign n34318 = ~n27206 ;
  assign n27210 = n34318 & n27208 ;
  assign n27211 = n27209 | n27210 ;
  assign n34319 = ~n27139 ;
  assign n27212 = n34319 & n27144 ;
  assign n27213 = n27211 | n27212 ;
  assign n27214 = n27211 & n27212 ;
  assign n34320 = ~n27214 ;
  assign n245 = n27213 & n34320 ;
  assign n34321 = ~n27210 ;
  assign n27216 = n34321 & n27213 ;
  assign n34322 = ~n27193 ;
  assign n27204 = n34322 & n27202 ;
  assign n27217 = n27201 | n27204 ;
  assign n34323 = ~n27180 ;
  assign n27218 = n27147 & n34323 ;
  assign n34324 = ~n27183 ;
  assign n27219 = n34324 & n27190 ;
  assign n27220 = n27218 | n27219 ;
  assign n5635 = n1457 & n5629 ;
  assign n1375 = x[125] & n1319 ;
  assign n1446 = x[126] & n1384 ;
  assign n27221 = n1375 | n1446 ;
  assign n27222 = x[127] & n1315 ;
  assign n27223 = n27221 | n27222 ;
  assign n27224 = n5635 | n27223 ;
  assign n34325 = ~n27224 ;
  assign n27225 = x[56] & n34325 ;
  assign n27226 = n30379 & n27224 ;
  assign n27227 = n27225 | n27226 ;
  assign n27228 = n27220 | n27227 ;
  assign n27229 = n27220 & n27227 ;
  assign n34326 = ~n27229 ;
  assign n27230 = n27228 & n34326 ;
  assign n27231 = n27169 | n27179 ;
  assign n5851 = n1217 & n5838 ;
  assign n1093 = x[122] & n1079 ;
  assign n1203 = x[123] & n1144 ;
  assign n27232 = n1093 | n1203 ;
  assign n27233 = x[124] & n1075 ;
  assign n27234 = n27232 | n27233 ;
  assign n27235 = n5851 | n27234 ;
  assign n34327 = ~n27235 ;
  assign n27236 = x[59] & n34327 ;
  assign n27237 = n30638 & n27235 ;
  assign n27238 = n27236 | n27237 ;
  assign n27152 = x[53] | n27151 ;
  assign n27239 = x[53] & n27151 ;
  assign n34328 = ~n27239 ;
  assign n27240 = n27152 & n34328 ;
  assign n308 = x[117] & n27215 ;
  assign n807 = x[118] & n805 ;
  assign n27241 = n308 | n807 ;
  assign n34329 = ~n27241 ;
  assign n27242 = n27240 & n34329 ;
  assign n34330 = ~n27240 ;
  assign n27243 = n34330 & n27241 ;
  assign n27244 = n27242 | n27243 ;
  assign n4998 = n1006 & n4985 ;
  assign n933 = x[119] & n900 ;
  assign n953 = x[120] & n949 ;
  assign n27245 = n933 | n953 ;
  assign n27246 = x[121] & n881 ;
  assign n27247 = n27245 | n27246 ;
  assign n27248 = n4998 | n27247 ;
  assign n34331 = ~n27248 ;
  assign n27249 = x[62] & n34331 ;
  assign n27250 = n30886 & n27248 ;
  assign n27251 = n27249 | n27250 ;
  assign n27252 = n27244 | n27251 ;
  assign n27253 = n27244 & n27251 ;
  assign n34332 = ~n27253 ;
  assign n27254 = n27252 & n34332 ;
  assign n27255 = n27158 & n27254 ;
  assign n27256 = n27158 | n27254 ;
  assign n34333 = ~n27255 ;
  assign n27257 = n34333 & n27256 ;
  assign n27258 = n27238 | n27257 ;
  assign n27259 = n27238 & n27257 ;
  assign n34334 = ~n27259 ;
  assign n27260 = n27258 & n34334 ;
  assign n34335 = ~n27231 ;
  assign n27261 = n34335 & n27260 ;
  assign n34336 = ~n27260 ;
  assign n27262 = n27231 & n34336 ;
  assign n27263 = n27261 | n27262 ;
  assign n27265 = n27230 & n27263 ;
  assign n27266 = n27230 | n27263 ;
  assign n34337 = ~n27265 ;
  assign n27267 = n34337 & n27266 ;
  assign n34338 = ~n27217 ;
  assign n27268 = n34338 & n27267 ;
  assign n34339 = ~n27267 ;
  assign n27269 = n27217 & n34339 ;
  assign n27270 = n27268 | n27269 ;
  assign n27271 = n27216 & n27270 ;
  assign n27272 = n27216 | n27270 ;
  assign n34340 = ~n27271 ;
  assign n246 = n34340 & n27272 ;
  assign n34341 = ~n27257 ;
  assign n27274 = n27238 & n34341 ;
  assign n27275 = n27262 | n27274 ;
  assign n1224 = n642 & n1217 ;
  assign n1130 = x[123] & n1079 ;
  assign n1204 = x[124] & n1144 ;
  assign n27276 = n1130 | n1204 ;
  assign n27277 = x[125] & n1075 ;
  assign n27278 = n27276 | n27277 ;
  assign n27279 = n1224 | n27278 ;
  assign n34342 = ~n27279 ;
  assign n27280 = x[59] & n34342 ;
  assign n27281 = n30638 & n27279 ;
  assign n27282 = n27280 | n27281 ;
  assign n34343 = ~n27244 ;
  assign n27283 = n34343 & n27251 ;
  assign n34344 = ~n27254 ;
  assign n27284 = n27158 & n34344 ;
  assign n27285 = n27283 | n27284 ;
  assign n309 = x[118] & n27215 ;
  assign n862 = x[119] & n805 ;
  assign n27286 = n309 | n862 ;
  assign n27287 = n30125 & n27151 ;
  assign n27288 = n27243 | n27287 ;
  assign n34345 = ~n27288 ;
  assign n27289 = n27286 & n34345 ;
  assign n34346 = ~n27286 ;
  assign n27290 = n34346 & n27288 ;
  assign n27291 = n27289 | n27290 ;
  assign n895 = x[122] & n881 ;
  assign n27292 = x[120] & n900 ;
  assign n27293 = x[121] & n949 ;
  assign n27294 = n27292 | n27293 ;
  assign n27295 = n895 | n27294 ;
  assign n27296 = n1006 & n5022 ;
  assign n27297 = n27295 | n27296 ;
  assign n27298 = n30886 & n27297 ;
  assign n34347 = ~n27297 ;
  assign n27299 = x[62] & n34347 ;
  assign n27300 = n27298 | n27299 ;
  assign n27301 = n27291 | n27300 ;
  assign n27302 = n27291 & n27300 ;
  assign n34348 = ~n27302 ;
  assign n27303 = n27301 & n34348 ;
  assign n27304 = n27285 | n27303 ;
  assign n27305 = n27285 & n27303 ;
  assign n34349 = ~n27305 ;
  assign n27306 = n27304 & n34349 ;
  assign n34350 = ~n27306 ;
  assign n27307 = n27282 & n34350 ;
  assign n34351 = ~n27282 ;
  assign n27308 = n34351 & n27304 ;
  assign n27309 = n34349 & n27308 ;
  assign n27310 = n27307 | n27309 ;
  assign n27311 = n27275 | n27310 ;
  assign n27312 = n27275 & n27310 ;
  assign n34352 = ~n27312 ;
  assign n27313 = n27311 & n34352 ;
  assign n6198 = n1457 & n6186 ;
  assign n1369 = x[126] & n1319 ;
  assign n27314 = x[127] & n1384 ;
  assign n27315 = n1369 | n27314 ;
  assign n27316 = n6198 | n27315 ;
  assign n34353 = ~n27316 ;
  assign n27317 = x[56] & n34353 ;
  assign n27318 = n30379 & n27316 ;
  assign n27319 = n27317 | n27318 ;
  assign n27320 = n27313 | n27319 ;
  assign n27321 = n27313 & n27319 ;
  assign n34354 = ~n27321 ;
  assign n27322 = n27320 & n34354 ;
  assign n34355 = ~n27263 ;
  assign n27264 = n27230 & n34355 ;
  assign n27323 = n27229 | n27264 ;
  assign n34356 = ~n27323 ;
  assign n27324 = n27322 & n34356 ;
  assign n34357 = ~n27322 ;
  assign n27325 = n34357 & n27323 ;
  assign n27326 = n27324 | n27325 ;
  assign n34358 = ~n27269 ;
  assign n27327 = n34358 & n27272 ;
  assign n27328 = n27326 | n27327 ;
  assign n27329 = n27326 & n27327 ;
  assign n34359 = ~n27329 ;
  assign n247 = n27328 & n34359 ;
  assign n5425 = n1006 & n5417 ;
  assign n934 = x[121] & n900 ;
  assign n968 = x[122] & n949 ;
  assign n27331 = n934 | n968 ;
  assign n27332 = x[123] & n881 ;
  assign n27333 = n27331 | n27332 ;
  assign n27334 = n5425 | n27333 ;
  assign n27335 = x[62] | n27334 ;
  assign n27336 = x[62] & n27334 ;
  assign n34360 = ~n27336 ;
  assign n27337 = n27335 & n34360 ;
  assign n310 = x[119] & n27215 ;
  assign n859 = x[120] & n805 ;
  assign n27338 = n310 | n859 ;
  assign n27339 = n27286 | n27338 ;
  assign n27340 = n27286 & n27338 ;
  assign n34361 = ~n27340 ;
  assign n27341 = n27339 & n34361 ;
  assign n27342 = n27337 & n27341 ;
  assign n27343 = n27337 | n27341 ;
  assign n34362 = ~n27342 ;
  assign n27344 = n34362 & n27343 ;
  assign n34363 = ~n27291 ;
  assign n27345 = n34363 & n27300 ;
  assign n27346 = n27290 | n27345 ;
  assign n34364 = ~n27346 ;
  assign n27347 = n27344 & n34364 ;
  assign n34365 = ~n27344 ;
  assign n27348 = n34365 & n27346 ;
  assign n27349 = n27347 | n27348 ;
  assign n5402 = n1217 & n5388 ;
  assign n1107 = x[124] & n1079 ;
  assign n1205 = x[125] & n1144 ;
  assign n27350 = n1107 | n1205 ;
  assign n27351 = x[126] & n1075 ;
  assign n27352 = n27350 | n27351 ;
  assign n27353 = n5402 | n27352 ;
  assign n34366 = ~n27353 ;
  assign n27354 = x[59] & n34366 ;
  assign n27355 = n30638 & n27353 ;
  assign n27356 = n27354 | n27355 ;
  assign n27357 = n27349 | n27356 ;
  assign n27358 = n27349 & n27356 ;
  assign n34367 = ~n27358 ;
  assign n27359 = n27357 & n34367 ;
  assign n34368 = ~n27303 ;
  assign n27360 = n27285 & n34368 ;
  assign n27361 = n27307 | n27360 ;
  assign n1383 = x[127] & n1319 ;
  assign n5373 = n1457 & n5360 ;
  assign n27362 = n1383 | n5373 ;
  assign n34369 = ~n27362 ;
  assign n27363 = x[56] & n34369 ;
  assign n27364 = n30379 & n27362 ;
  assign n27365 = n27363 | n27364 ;
  assign n27366 = n27361 | n27365 ;
  assign n27367 = n27361 & n27365 ;
  assign n34370 = ~n27367 ;
  assign n27368 = n27366 & n34370 ;
  assign n34371 = ~n27359 ;
  assign n27369 = n34371 & n27368 ;
  assign n34372 = ~n27368 ;
  assign n27370 = n27359 & n34372 ;
  assign n27371 = n27369 | n27370 ;
  assign n34373 = ~n27310 ;
  assign n27372 = n27275 & n34373 ;
  assign n34374 = ~n27313 ;
  assign n27373 = n34374 & n27319 ;
  assign n27374 = n27372 | n27373 ;
  assign n34375 = ~n27374 ;
  assign n27375 = n27371 & n34375 ;
  assign n34376 = ~n27371 ;
  assign n27376 = n34376 & n27374 ;
  assign n27377 = n27375 | n27376 ;
  assign n34377 = ~n27325 ;
  assign n27378 = n34377 & n27328 ;
  assign n27379 = n27377 & n27378 ;
  assign n27380 = n27377 | n27378 ;
  assign n34378 = ~n27379 ;
  assign n248 = n34378 & n27380 ;
  assign n34379 = ~n27349 ;
  assign n27404 = n34379 & n27356 ;
  assign n27405 = n27348 | n27404 ;
  assign n5632 = n1217 & n5629 ;
  assign n1143 = x[125] & n1079 ;
  assign n1206 = x[126] & n1144 ;
  assign n27406 = n1143 | n1206 ;
  assign n27407 = x[127] & n1075 ;
  assign n27408 = n27406 | n27407 ;
  assign n27409 = n5632 | n27408 ;
  assign n34380 = ~n27409 ;
  assign n27410 = x[59] & n34380 ;
  assign n27411 = n30638 & n27409 ;
  assign n27412 = n27410 | n27411 ;
  assign n27413 = n27405 | n27412 ;
  assign n27414 = n27405 & n27412 ;
  assign n34381 = ~n27414 ;
  assign n27415 = n27413 & n34381 ;
  assign n311 = x[120] & n27215 ;
  assign n809 = x[121] & n805 ;
  assign n27382 = n311 | n809 ;
  assign n27383 = x[56] | n27382 ;
  assign n27384 = x[56] & n27382 ;
  assign n34382 = ~n27384 ;
  assign n27385 = n27383 & n34382 ;
  assign n27386 = n27286 & n27385 ;
  assign n27387 = n27286 | n27385 ;
  assign n34383 = ~n27386 ;
  assign n27388 = n34383 & n27387 ;
  assign n27389 = n34346 & n27338 ;
  assign n34384 = ~n27341 ;
  assign n27390 = n27337 & n34384 ;
  assign n27391 = n27389 | n27390 ;
  assign n27392 = n27388 | n27391 ;
  assign n27393 = n27388 & n27391 ;
  assign n34385 = ~n27393 ;
  assign n27394 = n27392 & n34385 ;
  assign n5852 = n1006 & n5838 ;
  assign n947 = x[122] & n900 ;
  assign n969 = x[123] & n949 ;
  assign n27395 = n947 | n969 ;
  assign n27396 = x[124] & n881 ;
  assign n27397 = n27395 | n27396 ;
  assign n27398 = n5852 | n27397 ;
  assign n34386 = ~n27398 ;
  assign n27399 = x[62] & n34386 ;
  assign n27400 = n30886 & n27398 ;
  assign n27401 = n27399 | n27400 ;
  assign n34387 = ~n27394 ;
  assign n27403 = n34387 & n27401 ;
  assign n34388 = ~n27401 ;
  assign n27402 = n27394 & n34388 ;
  assign n34389 = ~n27402 ;
  assign n27416 = n34389 & n27415 ;
  assign n34390 = ~n27403 ;
  assign n27417 = n34390 & n27416 ;
  assign n34391 = ~n27417 ;
  assign n27418 = n27415 & n34391 ;
  assign n27419 = n27402 | n27417 ;
  assign n27420 = n27403 | n27419 ;
  assign n34392 = ~n27418 ;
  assign n27421 = n34392 & n27420 ;
  assign n27422 = n27367 | n27369 ;
  assign n34393 = ~n27422 ;
  assign n27423 = n27421 & n34393 ;
  assign n34394 = ~n27421 ;
  assign n27424 = n34394 & n27422 ;
  assign n27425 = n27423 | n27424 ;
  assign n34395 = ~n27376 ;
  assign n27426 = n34395 & n27380 ;
  assign n27427 = n27425 | n27426 ;
  assign n27428 = n27425 & n27426 ;
  assign n34396 = ~n27428 ;
  assign n249 = n27427 & n34396 ;
  assign n34397 = ~n27388 ;
  assign n27430 = n34397 & n27391 ;
  assign n27431 = n27403 | n27430 ;
  assign n312 = x[121] & n27215 ;
  assign n850 = x[122] & n805 ;
  assign n27432 = n312 | n850 ;
  assign n27433 = n30379 & n27382 ;
  assign n34398 = ~n27385 ;
  assign n27434 = n27286 & n34398 ;
  assign n27435 = n27433 | n27434 ;
  assign n27436 = n27432 | n27435 ;
  assign n27437 = n27432 & n27435 ;
  assign n34399 = ~n27437 ;
  assign n27438 = n27436 & n34399 ;
  assign n896 = x[125] & n881 ;
  assign n27439 = x[123] & n900 ;
  assign n27440 = x[124] & n949 ;
  assign n27441 = n27439 | n27440 ;
  assign n27442 = n896 | n27441 ;
  assign n27443 = n642 & n1006 ;
  assign n27444 = n27442 | n27443 ;
  assign n27445 = n30886 & n27444 ;
  assign n34400 = ~n27444 ;
  assign n27446 = x[62] & n34400 ;
  assign n27447 = n27445 | n27446 ;
  assign n27448 = n27438 | n27447 ;
  assign n27449 = n27438 & n27447 ;
  assign n34401 = ~n27449 ;
  assign n27450 = n27448 & n34401 ;
  assign n27451 = n27431 | n27450 ;
  assign n27452 = n27431 & n27450 ;
  assign n34402 = ~n27452 ;
  assign n27453 = n27451 & n34402 ;
  assign n6199 = n1217 & n6186 ;
  assign n1099 = x[126] & n1079 ;
  assign n27454 = x[127] & n1144 ;
  assign n27455 = n1099 | n27454 ;
  assign n27456 = n6199 | n27455 ;
  assign n34403 = ~n27456 ;
  assign n27457 = x[59] & n34403 ;
  assign n27458 = n30638 & n27456 ;
  assign n27459 = n27457 | n27458 ;
  assign n27460 = n27453 | n27459 ;
  assign n27461 = n27453 & n27459 ;
  assign n34404 = ~n27461 ;
  assign n27462 = n27460 & n34404 ;
  assign n27463 = n27414 | n27417 ;
  assign n34405 = ~n27463 ;
  assign n27464 = n27462 & n34405 ;
  assign n34406 = ~n27462 ;
  assign n27465 = n34406 & n27463 ;
  assign n27466 = n27464 | n27465 ;
  assign n34407 = ~n27424 ;
  assign n27467 = n34407 & n27427 ;
  assign n27468 = n27466 & n27467 ;
  assign n27469 = n27466 | n27467 ;
  assign n34408 = ~n27468 ;
  assign n250 = n34408 & n27469 ;
  assign n34409 = ~n27465 ;
  assign n27506 = n34409 & n27469 ;
  assign n34410 = ~n27450 ;
  assign n27471 = n27431 & n34410 ;
  assign n34411 = ~n27453 ;
  assign n27472 = n34411 & n27459 ;
  assign n27473 = n27471 | n27472 ;
  assign n34412 = ~n27432 ;
  assign n27477 = n34412 & n27435 ;
  assign n34413 = ~n27438 ;
  assign n27478 = n34413 & n27447 ;
  assign n27480 = n27477 | n27478 ;
  assign n313 = x[122] & n27215 ;
  assign n812 = x[123] & n805 ;
  assign n27474 = n313 | n812 ;
  assign n27476 = n34412 & n27474 ;
  assign n34414 = ~n27474 ;
  assign n27479 = n27432 & n34414 ;
  assign n27481 = n27476 | n27479 ;
  assign n27482 = n27480 & n27481 ;
  assign n34415 = ~n27476 ;
  assign n27483 = n34415 & n27480 ;
  assign n27484 = n27479 | n27483 ;
  assign n27485 = n27476 | n27484 ;
  assign n34416 = ~n27482 ;
  assign n27486 = n34416 & n27485 ;
  assign n5398 = n1006 & n5388 ;
  assign n910 = x[124] & n900 ;
  assign n976 = x[125] & n949 ;
  assign n27487 = n910 | n976 ;
  assign n27488 = x[126] & n881 ;
  assign n27489 = n27487 | n27488 ;
  assign n27490 = n5398 | n27489 ;
  assign n34417 = ~n27490 ;
  assign n27491 = x[62] & n34417 ;
  assign n27492 = n30886 & n27490 ;
  assign n27493 = n27491 | n27492 ;
  assign n1128 = x[127] & n1079 ;
  assign n5364 = n1217 & n5360 ;
  assign n27494 = n1128 | n5364 ;
  assign n34418 = ~n27494 ;
  assign n27495 = x[59] & n34418 ;
  assign n27496 = n30638 & n27494 ;
  assign n27497 = n27495 | n27496 ;
  assign n34419 = ~n27497 ;
  assign n27498 = n27493 & n34419 ;
  assign n34420 = ~n27493 ;
  assign n27499 = n34420 & n27497 ;
  assign n27500 = n27498 | n27499 ;
  assign n27502 = n27486 | n27500 ;
  assign n27503 = n27486 & n27500 ;
  assign n34421 = ~n27503 ;
  assign n27504 = n27502 & n34421 ;
  assign n27505 = n27473 & n27504 ;
  assign n27507 = n27473 | n27504 ;
  assign n34422 = ~n27505 ;
  assign n27508 = n34422 & n27507 ;
  assign n27509 = n27506 | n27508 ;
  assign n27510 = n27506 & n27507 ;
  assign n27511 = n34422 & n27510 ;
  assign n34423 = ~n27511 ;
  assign n251 = n27509 & n34423 ;
  assign n34424 = ~n27486 ;
  assign n27501 = n34424 & n27500 ;
  assign n27513 = n27493 & n27497 ;
  assign n27514 = n27501 | n27513 ;
  assign n27475 = x[59] | n27474 ;
  assign n27515 = x[59] & n27474 ;
  assign n34425 = ~n27515 ;
  assign n27516 = n27475 & n34425 ;
  assign n314 = x[123] & n27215 ;
  assign n824 = x[124] & n805 ;
  assign n27517 = n314 | n824 ;
  assign n34426 = ~n27517 ;
  assign n27518 = n27516 & n34426 ;
  assign n34427 = ~n27516 ;
  assign n27519 = n34427 & n27517 ;
  assign n27520 = n27518 | n27519 ;
  assign n5636 = n1006 & n5629 ;
  assign n944 = x[125] & n900 ;
  assign n996 = x[126] & n949 ;
  assign n27521 = n944 | n996 ;
  assign n27522 = x[127] & n881 ;
  assign n27523 = n27521 | n27522 ;
  assign n27524 = n5636 | n27523 ;
  assign n34428 = ~n27524 ;
  assign n27525 = x[62] & n34428 ;
  assign n27526 = n30886 & n27524 ;
  assign n27527 = n27525 | n27526 ;
  assign n27528 = n27520 | n27527 ;
  assign n27529 = n27520 & n27527 ;
  assign n34429 = ~n27529 ;
  assign n27530 = n27528 & n34429 ;
  assign n27531 = n27484 & n27530 ;
  assign n27532 = n27484 | n27530 ;
  assign n34430 = ~n27531 ;
  assign n27533 = n34430 & n27532 ;
  assign n27534 = n27514 & n27533 ;
  assign n34431 = ~n27504 ;
  assign n27535 = n27473 & n34431 ;
  assign n34432 = ~n27535 ;
  assign n27536 = n27509 & n34432 ;
  assign n27537 = n27514 | n27533 ;
  assign n27539 = n27536 & n27537 ;
  assign n34433 = ~n27534 ;
  assign n27540 = n34433 & n27539 ;
  assign n27538 = n34433 & n27537 ;
  assign n27541 = n27536 | n27538 ;
  assign n34434 = ~n27540 ;
  assign n252 = n34434 & n27541 ;
  assign n34435 = ~n27533 ;
  assign n27543 = n27514 & n34435 ;
  assign n34436 = ~n27543 ;
  assign n27544 = n27541 & n34436 ;
  assign n34437 = ~n27520 ;
  assign n27545 = n34437 & n27527 ;
  assign n34438 = ~n27530 ;
  assign n27546 = n27484 & n34438 ;
  assign n27547 = n27545 | n27546 ;
  assign n315 = x[124] & n27215 ;
  assign n806 = x[125] & n805 ;
  assign n27548 = n315 | n806 ;
  assign n27549 = n30638 & n27474 ;
  assign n27550 = n27519 | n27549 ;
  assign n34439 = ~n27550 ;
  assign n27551 = n27548 & n34439 ;
  assign n34440 = ~n27548 ;
  assign n27552 = n34440 & n27550 ;
  assign n27553 = n27551 | n27552 ;
  assign n6200 = n1006 & n6186 ;
  assign n27554 = x[126] & n900 ;
  assign n27555 = x[127] & n949 ;
  assign n27556 = n27554 | n27555 ;
  assign n27557 = n6200 | n27556 ;
  assign n34441 = ~n27557 ;
  assign n27558 = x[62] & n34441 ;
  assign n27559 = n30886 & n27557 ;
  assign n27560 = n27558 | n27559 ;
  assign n27561 = n27553 | n27560 ;
  assign n27562 = n27553 & n27560 ;
  assign n34442 = ~n27562 ;
  assign n27563 = n27561 & n34442 ;
  assign n27564 = n27547 & n27563 ;
  assign n27565 = n27547 | n27563 ;
  assign n34443 = ~n27564 ;
  assign n27566 = n34443 & n27565 ;
  assign n27567 = n27544 | n27566 ;
  assign n27568 = n27544 & n27565 ;
  assign n27569 = n34443 & n27568 ;
  assign n34444 = ~n27569 ;
  assign n253 = n27567 & n34444 ;
  assign n34445 = ~n27563 ;
  assign n27585 = n27547 & n34445 ;
  assign n34446 = ~n27585 ;
  assign n27586 = n27567 & n34446 ;
  assign n34447 = ~n27553 ;
  assign n27571 = n34447 & n27560 ;
  assign n27572 = n27552 | n27571 ;
  assign n316 = x[125] & n27215 ;
  assign n865 = x[126] & n805 ;
  assign n27573 = n316 | n865 ;
  assign n27574 = n27548 | n27573 ;
  assign n27575 = n27548 & n27573 ;
  assign n34448 = ~n27575 ;
  assign n27576 = n27574 & n34448 ;
  assign n948 = x[127] & n900 ;
  assign n5374 = n1006 & n5360 ;
  assign n27577 = n948 | n5374 ;
  assign n34449 = ~n27577 ;
  assign n27578 = x[62] & n34449 ;
  assign n27579 = n30886 & n27577 ;
  assign n27580 = n27578 | n27579 ;
  assign n34450 = ~n27580 ;
  assign n27581 = n27576 & n34450 ;
  assign n34451 = ~n27576 ;
  assign n27582 = n34451 & n27580 ;
  assign n27583 = n27581 | n27582 ;
  assign n27584 = n27572 & n27583 ;
  assign n27587 = n27572 | n27583 ;
  assign n34452 = ~n27584 ;
  assign n27588 = n34452 & n27587 ;
  assign n27589 = n27586 | n27588 ;
  assign n27590 = n27586 & n27587 ;
  assign n27591 = n34452 & n27590 ;
  assign n34453 = ~n27591 ;
  assign n254 = n27589 & n34453 ;
  assign n34454 = ~n27583 ;
  assign n27593 = n27572 & n34454 ;
  assign n34455 = ~n27593 ;
  assign n27594 = n27589 & n34455 ;
  assign n27595 = n34440 & n27573 ;
  assign n27596 = n27582 | n27595 ;
  assign n317 = x[126] & n27215 ;
  assign n866 = x[127] & n805 ;
  assign n27597 = n317 | n866 ;
  assign n34456 = ~n27597 ;
  assign n27598 = x[62] & n34456 ;
  assign n27599 = n30886 & n27597 ;
  assign n27600 = n27598 | n27599 ;
  assign n34457 = ~n27600 ;
  assign n27601 = n27548 & n34457 ;
  assign n27602 = n34440 & n27600 ;
  assign n27603 = n27601 | n27602 ;
  assign n34458 = ~n27603 ;
  assign n27604 = n27596 & n34458 ;
  assign n34459 = ~n27596 ;
  assign n27605 = n34459 & n27603 ;
  assign n27606 = n27604 | n27605 ;
  assign n27607 = n27594 | n27606 ;
  assign n27608 = n27594 & n27606 ;
  assign n34460 = ~n27608 ;
  assign n255 = n27607 & n34460 ;
  assign n27610 = n27599 | n27601 ;
  assign n27611 = x[127] & n27215 ;
  assign n27612 = n27610 & n27611 ;
  assign n27613 = n27610 | n27611 ;
  assign n34461 = ~n27612 ;
  assign n27614 = n34461 & n27613 ;
  assign n34462 = ~n27604 ;
  assign n27615 = n34462 & n27607 ;
  assign n27616 = n27614 & n27615 ;
  assign n27617 = n27614 | n27615 ;
  assign n34463 = ~n27616 ;
  assign n256 = n34463 & n27617 ;
  assign y[0] = n129 ;
  assign y[1] = n130 ;
  assign y[2] = n131 ;
  assign y[3] = n132 ;
  assign y[4] = n133 ;
  assign y[5] = n134 ;
  assign y[6] = n135 ;
  assign y[7] = n136 ;
  assign y[8] = n137 ;
  assign y[9] = n138 ;
  assign y[10] = n139 ;
  assign y[11] = n140 ;
  assign y[12] = n141 ;
  assign y[13] = n142 ;
  assign y[14] = n143 ;
  assign y[15] = n144 ;
  assign y[16] = n145 ;
  assign y[17] = n146 ;
  assign y[18] = n147 ;
  assign y[19] = n148 ;
  assign y[20] = n149 ;
  assign y[21] = n150 ;
  assign y[22] = n151 ;
  assign y[23] = n152 ;
  assign y[24] = n153 ;
  assign y[25] = n154 ;
  assign y[26] = n155 ;
  assign y[27] = n156 ;
  assign y[28] = n157 ;
  assign y[29] = n158 ;
  assign y[30] = n159 ;
  assign y[31] = n160 ;
  assign y[32] = n161 ;
  assign y[33] = n162 ;
  assign y[34] = n163 ;
  assign y[35] = n164 ;
  assign y[36] = n165 ;
  assign y[37] = n166 ;
  assign y[38] = n167 ;
  assign y[39] = n168 ;
  assign y[40] = n169 ;
  assign y[41] = n170 ;
  assign y[42] = n171 ;
  assign y[43] = n172 ;
  assign y[44] = n173 ;
  assign y[45] = n174 ;
  assign y[46] = n175 ;
  assign y[47] = n176 ;
  assign y[48] = n177 ;
  assign y[49] = n178 ;
  assign y[50] = n179 ;
  assign y[51] = n180 ;
  assign y[52] = n181 ;
  assign y[53] = n182 ;
  assign y[54] = n183 ;
  assign y[55] = n184 ;
  assign y[56] = n185 ;
  assign y[57] = n186 ;
  assign y[58] = n187 ;
  assign y[59] = n188 ;
  assign y[60] = n189 ;
  assign y[61] = n190 ;
  assign y[62] = n191 ;
  assign y[63] = n192 ;
  assign y[64] = n193 ;
  assign y[65] = n194 ;
  assign y[66] = n195 ;
  assign y[67] = n196 ;
  assign y[68] = n197 ;
  assign y[69] = n198 ;
  assign y[70] = n199 ;
  assign y[71] = n200 ;
  assign y[72] = n201 ;
  assign y[73] = n202 ;
  assign y[74] = n203 ;
  assign y[75] = n204 ;
  assign y[76] = n205 ;
  assign y[77] = n206 ;
  assign y[78] = n207 ;
  assign y[79] = n208 ;
  assign y[80] = n209 ;
  assign y[81] = n210 ;
  assign y[82] = n211 ;
  assign y[83] = n212 ;
  assign y[84] = n213 ;
  assign y[85] = n214 ;
  assign y[86] = n215 ;
  assign y[87] = n216 ;
  assign y[88] = n217 ;
  assign y[89] = n218 ;
  assign y[90] = n219 ;
  assign y[91] = n220 ;
  assign y[92] = n221 ;
  assign y[93] = n222 ;
  assign y[94] = n223 ;
  assign y[95] = n224 ;
  assign y[96] = n225 ;
  assign y[97] = n226 ;
  assign y[98] = n227 ;
  assign y[99] = n228 ;
  assign y[100] = n229 ;
  assign y[101] = n230 ;
  assign y[102] = n231 ;
  assign y[103] = n232 ;
  assign y[104] = n233 ;
  assign y[105] = n234 ;
  assign y[106] = n235 ;
  assign y[107] = n236 ;
  assign y[108] = n237 ;
  assign y[109] = n238 ;
  assign y[110] = n239 ;
  assign y[111] = n240 ;
  assign y[112] = n241 ;
  assign y[113] = n242 ;
  assign y[114] = n243 ;
  assign y[115] = n244 ;
  assign y[116] = n245 ;
  assign y[117] = n246 ;
  assign y[118] = n247 ;
  assign y[119] = n248 ;
  assign y[120] = n249 ;
  assign y[121] = n250 ;
  assign y[122] = n251 ;
  assign y[123] = n252 ;
  assign y[124] = n253 ;
  assign y[125] = n254 ;
  assign y[126] = n255 ;
  assign y[127] = n256 ;
endmodule
