module sin( input [23:0] x , output [24:0] y );
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 ;
  assign n4081 = x[21] & x[22] ;
  assign n5243 = x[1] | x[2] ;
  assign n5294 = x[0] | n5243 ;
  assign n5333 = x[3] | n5294 ;
  assign n5378 = x[4] | n5333 ;
  assign n5401 = x[5] | n5378 ;
  assign n5440 = x[6] | n5401 ;
  assign n5454 = x[7] | n5440 ;
  assign n6771 = x[8] | n5454 ;
  assign n50 = x[9] | n6771 ;
  assign n52 = x[10] | n50 ;
  assign n53 = x[11] | n52 ;
  assign n55 = x[12] | n53 ;
  assign n56 = x[13] | n55 ;
  assign n58 = x[14] | n56 ;
  assign n60 = x[15] | n58 ;
  assign n61 = x[16] | n60 ;
  assign n62 = x[17] | n61 ;
  assign n64 = x[18] | n62 ;
  assign n65 = x[19] | n64 ;
  assign n67 = x[20] | n65 ;
  assign n5471 = ~n67 ;
  assign n68 = x[21] & n5471 ;
  assign n5472 = ~x[21] ;
  assign n70 = n5472 & n67 ;
  assign n71 = n68 | n70 ;
  assign n5473 = ~x[22] ;
  assign n72 = n5473 & n71 ;
  assign n73 = n4081 | n72 ;
  assign n4212 = x[20] & x[22] ;
  assign n5474 = ~n65 ;
  assign n66 = x[20] & n5474 ;
  assign n5475 = ~x[20] ;
  assign n74 = n5475 & n65 ;
  assign n75 = n66 | n74 ;
  assign n76 = n5473 & n75 ;
  assign n77 = n4212 | n76 ;
  assign n78 = n73 | n77 ;
  assign n4326 = x[15] & x[22] ;
  assign n59 = x[15] & n58 ;
  assign n79 = n5473 & n60 ;
  assign n5476 = ~n59 ;
  assign n81 = n5476 & n79 ;
  assign n82 = n4326 | n81 ;
  assign n83 = n78 | n82 ;
  assign n84 = n5473 & n64 ;
  assign n85 = x[19] & n84 ;
  assign n86 = x[19] | n84 ;
  assign n5477 = ~n85 ;
  assign n87 = n5477 & n86 ;
  assign n4423 = x[18] & x[22] ;
  assign n63 = x[18] & n62 ;
  assign n5478 = ~n63 ;
  assign n88 = n5478 & n84 ;
  assign n89 = n4423 | n88 ;
  assign n91 = n87 & n89 ;
  assign n92 = n5473 & n61 ;
  assign n93 = x[17] & n92 ;
  assign n94 = x[17] | n92 ;
  assign n5479 = ~n93 ;
  assign n95 = n5479 & n94 ;
  assign n80 = x[16] & n79 ;
  assign n96 = x[16] | n79 ;
  assign n5480 = ~n80 ;
  assign n97 = n5480 & n96 ;
  assign n5481 = ~n97 ;
  assign n99 = n95 & n5481 ;
  assign n100 = n91 & n99 ;
  assign n5482 = ~n83 ;
  assign n101 = n5482 & n100 ;
  assign n102 = n95 | n97 ;
  assign n5483 = ~n102 ;
  assign n103 = n91 & n5483 ;
  assign n4532 = n5475 & x[22] ;
  assign n104 = x[22] | n75 ;
  assign n5484 = ~n4532 ;
  assign n105 = n5484 & n104 ;
  assign n5485 = ~n73 ;
  assign n106 = n5485 & n105 ;
  assign n5486 = ~n82 ;
  assign n107 = n5486 & n106 ;
  assign n108 = n103 & n107 ;
  assign n5487 = ~n89 ;
  assign n90 = n87 & n5487 ;
  assign n109 = n90 & n5483 ;
  assign n110 = n107 & n109 ;
  assign n111 = n82 & n106 ;
  assign n5488 = ~n87 ;
  assign n112 = n5488 & n89 ;
  assign n113 = n5483 & n112 ;
  assign n114 = n111 & n113 ;
  assign n4638 = n5472 & x[22] ;
  assign n115 = x[22] | n71 ;
  assign n5489 = ~n4638 ;
  assign n116 = n5489 & n115 ;
  assign n5490 = ~n77 ;
  assign n117 = n5490 & n116 ;
  assign n118 = n82 & n117 ;
  assign n5491 = ~n95 ;
  assign n98 = n5491 & n97 ;
  assign n119 = n90 & n98 ;
  assign n120 = n118 & n119 ;
  assign n121 = n105 & n116 ;
  assign n122 = n82 & n121 ;
  assign n123 = n90 & n99 ;
  assign n124 = n122 & n123 ;
  assign n125 = n5486 & n121 ;
  assign n126 = n100 & n125 ;
  assign n5492 = ~n78 ;
  assign n127 = n5492 & n82 ;
  assign n128 = n99 & n112 ;
  assign n129 = n127 & n128 ;
  assign n130 = n100 & n118 ;
  assign n131 = n119 & n122 ;
  assign n132 = n95 & n97 ;
  assign n133 = n112 & n132 ;
  assign n134 = n122 & n133 ;
  assign n135 = n125 & n133 ;
  assign n136 = n119 & n125 ;
  assign n137 = n125 & n128 ;
  assign n138 = n136 | n137 ;
  assign n139 = n100 & n107 ;
  assign n140 = n91 & n98 ;
  assign n141 = n125 & n140 ;
  assign n142 = n139 | n141 ;
  assign n143 = n100 & n111 ;
  assign n144 = n98 & n112 ;
  assign n145 = n107 & n144 ;
  assign n146 = n143 | n145 ;
  assign n147 = n123 & n125 ;
  assign n148 = n90 & n132 ;
  assign n149 = n125 & n148 ;
  assign n150 = n147 | n149 ;
  assign n151 = n127 & n133 ;
  assign n152 = n100 & n122 ;
  assign n153 = n151 | n152 ;
  assign n154 = n150 | n153 ;
  assign n155 = n146 | n154 ;
  assign n156 = n142 | n155 ;
  assign n157 = n138 | n156 ;
  assign n158 = n135 | n157 ;
  assign n159 = n134 | n158 ;
  assign n160 = n131 | n159 ;
  assign n161 = n130 | n160 ;
  assign n162 = n129 | n161 ;
  assign n163 = n107 & n140 ;
  assign n164 = n118 & n148 ;
  assign n165 = n5482 & n148 ;
  assign n166 = n111 & n119 ;
  assign n167 = n87 | n89 ;
  assign n168 = n102 | n167 ;
  assign n5493 = ~n168 ;
  assign n169 = n111 & n5493 ;
  assign n170 = n5486 & n117 ;
  assign n171 = n148 & n170 ;
  assign n172 = n103 & n122 ;
  assign n173 = n122 & n140 ;
  assign n174 = n113 & n170 ;
  assign n175 = n103 & n125 ;
  assign n176 = n174 | n175 ;
  assign n177 = n173 | n176 ;
  assign n178 = n172 | n177 ;
  assign n179 = n171 | n178 ;
  assign n180 = n169 | n179 ;
  assign n181 = n166 | n180 ;
  assign n182 = n165 | n181 ;
  assign n183 = n103 & n118 ;
  assign n5494 = ~n167 ;
  assign n184 = n132 & n5494 ;
  assign n186 = n125 & n184 ;
  assign n187 = n183 | n186 ;
  assign n188 = n107 & n148 ;
  assign n189 = n113 & n118 ;
  assign n190 = n118 & n123 ;
  assign n191 = n98 & n5494 ;
  assign n192 = n122 & n191 ;
  assign n193 = n91 & n132 ;
  assign n194 = n125 & n193 ;
  assign n195 = n192 | n194 ;
  assign n196 = n190 | n195 ;
  assign n197 = n189 | n196 ;
  assign n198 = n188 | n197 ;
  assign n199 = n187 | n198 ;
  assign n200 = n182 | n199 ;
  assign n201 = n164 | n200 ;
  assign n202 = n163 | n201 ;
  assign n203 = n99 & n5494 ;
  assign n204 = n111 & n203 ;
  assign n205 = n118 & n128 ;
  assign n206 = n125 & n144 ;
  assign n207 = n205 | n206 ;
  assign n208 = n204 | n207 ;
  assign n209 = n127 & n144 ;
  assign n210 = n111 & n193 ;
  assign n211 = n5493 & n170 ;
  assign n212 = n122 & n5493 ;
  assign n213 = n113 & n127 ;
  assign n214 = n107 & n123 ;
  assign n215 = n118 & n144 ;
  assign n216 = n103 & n170 ;
  assign n217 = n122 & n184 ;
  assign n218 = n122 & n128 ;
  assign n219 = n122 & n144 ;
  assign n220 = n125 & n191 ;
  assign n221 = n119 & n127 ;
  assign n222 = n111 & n123 ;
  assign n223 = n118 & n140 ;
  assign n224 = n100 & n170 ;
  assign n225 = n122 & n148 ;
  assign n226 = n109 & n122 ;
  assign n227 = n225 | n226 ;
  assign n228 = n224 | n227 ;
  assign n229 = n223 | n228 ;
  assign n230 = n222 | n229 ;
  assign n231 = n221 | n230 ;
  assign n232 = n111 & n184 ;
  assign n233 = n100 & n127 ;
  assign n234 = n232 | n233 ;
  assign n235 = n127 & n184 ;
  assign n236 = n127 & n203 ;
  assign n237 = n235 | n236 ;
  assign n238 = n234 | n237 ;
  assign n239 = n231 | n238 ;
  assign n240 = n220 | n239 ;
  assign n241 = n219 | n240 ;
  assign n242 = n218 | n241 ;
  assign n243 = n217 | n242 ;
  assign n244 = n216 | n243 ;
  assign n245 = n215 | n244 ;
  assign n246 = n214 | n245 ;
  assign n247 = n213 | n246 ;
  assign n248 = n212 | n247 ;
  assign n249 = n211 | n248 ;
  assign n250 = n210 | n249 ;
  assign n251 = n209 | n250 ;
  assign n252 = n170 & n191 ;
  assign n253 = n118 & n193 ;
  assign n254 = n252 | n253 ;
  assign n255 = n109 & n170 ;
  assign n256 = n5482 & n191 ;
  assign n257 = n255 | n256 ;
  assign n258 = n254 | n257 ;
  assign n259 = n251 | n258 ;
  assign n260 = n208 | n259 ;
  assign n261 = n202 | n260 ;
  assign n262 = n162 | n261 ;
  assign n263 = n126 | n262 ;
  assign n264 = n124 | n263 ;
  assign n265 = n120 | n264 ;
  assign n266 = n114 | n265 ;
  assign n267 = n110 | n266 ;
  assign n268 = n108 | n267 ;
  assign n269 = n101 | n268 ;
  assign n270 = n5473 & n5378 ;
  assign n271 = x[5] & n270 ;
  assign n273 = x[5] | n270 ;
  assign n5495 = ~n271 ;
  assign n274 = n5495 & n273 ;
  assign n4731 = x[4] & x[22] ;
  assign n5355 = x[4] & n5333 ;
  assign n5496 = ~n5355 ;
  assign n272 = n5496 & n270 ;
  assign n275 = n4731 | n272 ;
  assign n279 = n5473 & n5294 ;
  assign n280 = x[3] & n279 ;
  assign n281 = x[3] | n279 ;
  assign n5497 = ~n280 ;
  assign n282 = n5497 & n281 ;
  assign n5498 = ~n275 ;
  assign n283 = n5498 & n282 ;
  assign n5499 = ~n282 ;
  assign n2559 = n275 & n5499 ;
  assign n2560 = n283 | n2559 ;
  assign n276 = n274 | n275 ;
  assign n277 = n274 & n275 ;
  assign n5500 = ~n277 ;
  assign n278 = n276 & n5500 ;
  assign n3924 = x[2] & x[22] ;
  assign n284 = x[0] | x[1] ;
  assign n285 = x[2] & n284 ;
  assign n5501 = ~n285 ;
  assign n286 = n279 & n5501 ;
  assign n287 = n3924 | n286 ;
  assign n5502 = ~n287 ;
  assign n288 = n282 & n5502 ;
  assign n290 = n5499 & n287 ;
  assign n291 = n288 | n290 ;
  assign n5503 = ~n291 ;
  assign n2561 = n278 & n5503 ;
  assign n5504 = ~n2560 ;
  assign n2562 = n5504 & n2561 ;
  assign n355 = n107 & n203 ;
  assign n294 = n103 & n111 ;
  assign n457 = n118 & n191 ;
  assign n468 = n123 & n127 ;
  assign n324 = n133 & n170 ;
  assign n414 = n140 & n170 ;
  assign n391 = n122 & n193 ;
  assign n405 = n113 & n125 ;
  assign n1006 = n220 | n405 ;
  assign n1007 = n391 | n1006 ;
  assign n1008 = n226 | n1007 ;
  assign n1009 = n414 | n1008 ;
  assign n332 = n107 & n191 ;
  assign n345 = n128 & n170 ;
  assign n494 = n111 & n191 ;
  assign n1137 = n345 | n494 ;
  assign n1138 = n332 | n1137 ;
  assign n552 = n5482 & n203 ;
  assign n445 = n118 & n5493 ;
  assign n1139 = n224 | n445 ;
  assign n1140 = n552 | n1139 ;
  assign n471 = n5482 & n140 ;
  assign n502 = n107 & n119 ;
  assign n340 = n170 & n184 ;
  assign n1141 = n172 | n340 ;
  assign n1142 = n502 | n1141 ;
  assign n1143 = n471 | n1142 ;
  assign n1144 = n1140 | n1143 ;
  assign n1145 = n1138 | n1144 ;
  assign n1146 = n1009 | n1145 ;
  assign n1147 = n146 | n1146 ;
  assign n1148 = n194 | n1147 ;
  assign n1149 = n324 | n1148 ;
  assign n1150 = n210 | n1149 ;
  assign n1151 = n468 | n1150 ;
  assign n553 = n5482 & n128 ;
  assign n505 = n107 & n128 ;
  assign n295 = n109 & n111 ;
  assign n370 = n101 | n213 ;
  assign n599 = n138 | n370 ;
  assign n600 = n218 | n599 ;
  assign n601 = n131 | n600 ;
  assign n602 = n169 | n601 ;
  assign n603 = n295 | n602 ;
  assign n604 = n505 | n603 ;
  assign n605 = n553 | n604 ;
  assign n354 = n107 & n133 ;
  assign n356 = n107 & n113 ;
  assign n347 = n123 & n170 ;
  assign n446 = n111 & n148 ;
  assign n357 = n118 & n184 ;
  assign n986 = n166 | n357 ;
  assign n987 = n446 | n986 ;
  assign n988 = n152 | n987 ;
  assign n989 = n347 | n988 ;
  assign n990 = n216 | n989 ;
  assign n991 = n232 | n990 ;
  assign n992 = n356 | n991 ;
  assign n993 = n354 | n992 ;
  assign n752 = n127 & n191 ;
  assign n753 = n120 | n164 ;
  assign n754 = n214 | n753 ;
  assign n755 = n752 | n754 ;
  assign n309 = n170 & n193 ;
  assign n412 = n125 & n5493 ;
  assign n636 = n309 | n412 ;
  assign n353 = n107 & n5493 ;
  assign n473 = n233 | n353 ;
  assign n314 = n122 & n203 ;
  assign n315 = n126 | n314 ;
  assign n316 = n205 | n315 ;
  assign n469 = n5482 & n103 ;
  assign n809 = n108 | n173 ;
  assign n810 = n469 | n809 ;
  assign n2214 = n142 | n810 ;
  assign n2215 = n316 | n2214 ;
  assign n2216 = n473 | n2215 ;
  assign n2217 = n636 | n2216 ;
  assign n2218 = n755 | n2217 ;
  assign n2219 = n993 | n2218 ;
  assign n2220 = n605 | n2219 ;
  assign n2221 = n1151 | n2220 ;
  assign n2222 = n457 | n2221 ;
  assign n2223 = n294 | n2222 ;
  assign n2224 = n355 | n2223 ;
  assign n2225 = n165 | n2224 ;
  assign n2226 = n235 | n2225 ;
  assign n668 = n5473 & n52 ;
  assign n669 = x[11] & n668 ;
  assign n671 = x[11] | n668 ;
  assign n5505 = ~n669 ;
  assign n672 = n5505 & n671 ;
  assign n444 = n5482 & n119 ;
  assign n365 = n5482 & n123 ;
  assign n447 = n188 | n446 ;
  assign n448 = n111 & n140 ;
  assign n449 = n294 | n448 ;
  assign n450 = n163 | n449 ;
  assign n451 = n447 | n450 ;
  assign n452 = n143 | n451 ;
  assign n453 = n252 | n340 ;
  assign n454 = n222 | n453 ;
  assign n455 = n210 | n454 ;
  assign n456 = n139 | n455 ;
  assign n297 = n118 & n203 ;
  assign n458 = n297 | n457 ;
  assign n344 = n107 & n193 ;
  assign n346 = n344 | n345 ;
  assign n367 = n170 & n203 ;
  assign n459 = n357 | n367 ;
  assign n460 = n346 | n459 ;
  assign n461 = n458 | n460 ;
  assign n462 = n456 | n461 ;
  assign n463 = n452 | n462 ;
  assign n464 = n211 | n463 ;
  assign n465 = n445 | n464 ;
  assign n466 = n108 | n465 ;
  assign n467 = n109 & n127 ;
  assign n293 = n127 & n148 ;
  assign n470 = n127 & n193 ;
  assign n364 = n5482 & n193 ;
  assign n326 = n144 & n170 ;
  assign n472 = n174 | n326 ;
  assign n474 = n189 | n215 ;
  assign n475 = n169 | n474 ;
  assign n339 = n103 & n127 ;
  assign n476 = n127 & n140 ;
  assign n477 = n339 | n476 ;
  assign n478 = n475 | n477 ;
  assign n479 = n473 | n478 ;
  assign n480 = n472 | n479 ;
  assign n481 = n101 | n480 ;
  assign n482 = n364 | n481 ;
  assign n483 = n471 | n482 ;
  assign n484 = n470 | n483 ;
  assign n485 = n469 | n484 ;
  assign n486 = n165 | n485 ;
  assign n487 = n293 | n486 ;
  assign n488 = n468 | n487 ;
  assign n489 = n467 | n488 ;
  assign n490 = n466 | n489 ;
  assign n491 = n365 | n490 ;
  assign n492 = n444 | n491 ;
  assign n493 = n221 | n492 ;
  assign n312 = n107 & n184 ;
  assign n495 = n114 | n332 ;
  assign n496 = n494 | n495 ;
  assign n497 = n355 | n496 ;
  assign n498 = n312 | n497 ;
  assign n499 = n232 | n498 ;
  assign n500 = n204 | n499 ;
  assign n501 = n356 | n500 ;
  assign n299 = n111 & n128 ;
  assign n503 = n111 & n133 ;
  assign n504 = n214 | n503 ;
  assign n358 = n111 & n144 ;
  assign n506 = n354 | n358 ;
  assign n507 = n505 | n506 ;
  assign n508 = n504 | n507 ;
  assign n509 = n299 | n508 ;
  assign n510 = n295 | n509 ;
  assign n511 = n166 | n510 ;
  assign n512 = n110 | n511 ;
  assign n513 = n502 | n512 ;
  assign n514 = n466 | n513 ;
  assign n515 = n474 | n514 ;
  assign n516 = n472 | n515 ;
  assign n517 = n501 | n516 ;
  assign n518 = n145 | n517 ;
  assign n5506 = ~n518 ;
  assign n519 = n493 & n5506 ;
  assign n5507 = ~n493 ;
  assign n537 = n5507 & n518 ;
  assign n538 = n519 | n537 ;
  assign n325 = n125 & n203 ;
  assign n392 = n190 | n347 ;
  assign n310 = n118 & n133 ;
  assign n311 = n219 | n310 ;
  assign n334 = n109 & n125 ;
  assign n393 = n171 | n334 ;
  assign n394 = n205 | n324 ;
  assign n395 = n393 | n394 ;
  assign n396 = n311 | n395 ;
  assign n397 = n138 | n396 ;
  assign n398 = n206 | n397 ;
  assign n399 = n226 | n398 ;
  assign n400 = n392 | n399 ;
  assign n401 = n164 | n400 ;
  assign n402 = n113 & n122 ;
  assign n333 = n109 & n118 ;
  assign n403 = n134 | n255 ;
  assign n404 = n333 | n403 ;
  assign n296 = n119 & n170 ;
  assign n406 = n135 | n405 ;
  assign n407 = n218 | n406 ;
  assign n408 = n296 | n407 ;
  assign n409 = n404 | n408 ;
  assign n410 = n402 | n409 ;
  assign n411 = n120 | n410 ;
  assign n413 = n253 | n412 ;
  assign n415 = n150 | n187 ;
  assign n416 = n124 | n415 ;
  assign n417 = n217 | n416 ;
  assign n418 = n223 | n417 ;
  assign n419 = n414 | n418 ;
  assign n420 = n216 | n419 ;
  assign n421 = n413 | n420 ;
  assign n422 = n411 | n421 ;
  assign n423 = n220 | n422 ;
  assign n424 = n141 | n423 ;
  assign n425 = n126 | n424 ;
  assign n426 = n173 | n425 ;
  assign n427 = n212 | n426 ;
  assign n428 = n131 | n427 ;
  assign n429 = n152 | n192 ;
  assign n430 = n175 | n225 ;
  assign n431 = n172 | n430 ;
  assign n432 = n309 | n431 ;
  assign n433 = n224 | n432 ;
  assign n434 = n130 | n433 ;
  assign n435 = n429 | n434 ;
  assign n436 = n428 | n435 ;
  assign n437 = n401 | n436 ;
  assign n438 = n325 | n437 ;
  assign n439 = n194 | n438 ;
  assign n440 = n314 | n439 ;
  assign n441 = n391 | n440 ;
  assign n541 = n493 | n518 ;
  assign n5508 = ~n441 ;
  assign n542 = n5508 & n541 ;
  assign n5509 = ~n542 ;
  assign n685 = n538 & n5509 ;
  assign n687 = n672 & n685 ;
  assign n520 = n493 & n518 ;
  assign n5510 = ~n520 ;
  assign n545 = n441 & n5510 ;
  assign n694 = n538 | n545 ;
  assign n4984 = x[10] & x[22] ;
  assign n51 = x[10] & n50 ;
  assign n5511 = ~n51 ;
  assign n670 = n5511 & n668 ;
  assign n859 = n4984 | n670 ;
  assign n5512 = ~n859 ;
  assign n863 = n694 & n5512 ;
  assign n543 = n538 | n542 ;
  assign n927 = n543 & n859 ;
  assign n928 = n863 | n927 ;
  assign n5513 = ~n545 ;
  assign n692 = n538 & n5513 ;
  assign n5514 = ~n672 ;
  assign n929 = n5514 & n692 ;
  assign n5515 = ~n929 ;
  assign n930 = n928 & n5515 ;
  assign n5516 = ~n687 ;
  assign n931 = n5516 & n930 ;
  assign n342 = n127 & n5493 ;
  assign n745 = n220 | n412 ;
  assign n746 = n217 | n745 ;
  assign n747 = n356 | n746 ;
  assign n748 = n163 | n747 ;
  assign n749 = n469 | n748 ;
  assign n750 = n365 | n749 ;
  assign n751 = n342 | n750 ;
  assign n348 = n5482 & n109 ;
  assign n756 = n334 | n494 ;
  assign n757 = n502 | n756 ;
  assign n758 = n505 | n757 ;
  assign n759 = n348 | n758 ;
  assign n760 = n233 | n759 ;
  assign n761 = n475 | n760 ;
  assign n762 = n755 | n761 ;
  assign n763 = n136 | n762 ;
  assign n764 = n503 | n763 ;
  assign n765 = n294 | n764 ;
  assign n766 = n204 | n765 ;
  assign n767 = n101 | n766 ;
  assign n768 = n236 | n767 ;
  assign n551 = n5482 & n133 ;
  assign n769 = n129 | n295 ;
  assign n644 = n135 | n226 ;
  assign n770 = n345 | n644 ;
  assign n771 = n347 | n770 ;
  assign n772 = n216 | n771 ;
  assign n773 = n145 | n772 ;
  assign n774 = n174 | n209 ;
  assign n775 = n213 | n774 ;
  assign n776 = n210 | n471 ;
  assign n777 = n775 | n776 ;
  assign n778 = n773 | n777 ;
  assign n779 = n769 | n778 ;
  assign n780 = n186 | n779 ;
  assign n781 = n255 | n780 ;
  assign n782 = n139 | n781 ;
  assign n783 = n551 | n782 ;
  assign n784 = n444 | n783 ;
  assign n785 = n134 | n310 ;
  assign n786 = n446 | n785 ;
  assign n787 = n312 | n786 ;
  assign n788 = n165 | n787 ;
  assign n789 = n470 | n788 ;
  assign n790 = n212 | n402 ;
  assign n791 = n299 | n790 ;
  assign n792 = n252 | n297 ;
  assign n793 = n223 | n792 ;
  assign n794 = n791 | n793 ;
  assign n795 = n789 | n794 ;
  assign n796 = n784 | n795 ;
  assign n797 = n768 | n796 ;
  assign n798 = n751 | n797 ;
  assign n799 = n405 | n798 ;
  assign n800 = n224 | n799 ;
  assign n801 = n130 | n800 ;
  assign n802 = n235 | n801 ;
  assign n932 = n163 | n445 ;
  assign n933 = n142 | n932 ;
  assign n934 = n551 | n933 ;
  assign n935 = n236 | n934 ;
  assign n936 = n293 | n935 ;
  assign n313 = n110 | n312 ;
  assign n317 = n313 | n316 ;
  assign n318 = n311 | n317 ;
  assign n319 = n309 | n318 ;
  assign n320 = n210 | n319 ;
  assign n300 = n108 | n299 ;
  assign n937 = n171 | n469 ;
  assign n938 = n220 | n937 ;
  assign n939 = n347 | n938 ;
  assign n940 = n342 | n939 ;
  assign n941 = n300 | n940 ;
  assign n942 = n320 | n941 ;
  assign n943 = n936 | n942 ;
  assign n944 = n149 | n943 ;
  assign n945 = n194 | n944 ;
  assign n946 = n183 | n945 ;
  assign n947 = n503 | n946 ;
  assign n948 = n494 | n947 ;
  assign n949 = n151 | n948 ;
  assign n950 = n367 | n467 ;
  assign n951 = n344 | n950 ;
  assign n952 = n444 | n951 ;
  assign n588 = n5482 & n184 ;
  assign n953 = n124 | n404 ;
  assign n954 = n214 | n953 ;
  assign n955 = n588 | n954 ;
  assign n956 = n364 | n955 ;
  assign n957 = n136 | n324 ;
  assign n560 = n232 | n470 ;
  assign n561 = n235 | n560 ;
  assign n637 = n173 | n502 ;
  assign n958 = n561 | n637 ;
  assign n959 = n957 | n958 ;
  assign n960 = n956 | n959 ;
  assign n961 = n952 | n960 ;
  assign n962 = n217 | n961 ;
  assign n963 = n296 | n962 ;
  assign n964 = n145 | n963 ;
  assign n965 = n174 | n212 ;
  assign n966 = n216 | n965 ;
  assign n967 = n190 | n966 ;
  assign n968 = n130 | n967 ;
  assign n969 = n752 | n968 ;
  assign n970 = n339 | n969 ;
  assign n321 = n83 | n168 ;
  assign n5517 = ~n120 ;
  assign n322 = n5517 & n321 ;
  assign n971 = n188 | n391 ;
  assign n972 = n233 | n971 ;
  assign n973 = n152 | n402 ;
  assign n974 = n348 | n973 ;
  assign n571 = n164 | n218 ;
  assign n572 = n189 | n571 ;
  assign n975 = n495 | n572 ;
  assign n976 = n974 | n975 ;
  assign n977 = n972 | n976 ;
  assign n5518 = ~n977 ;
  assign n978 = n322 & n5518 ;
  assign n5519 = ~n970 ;
  assign n979 = n5519 & n978 ;
  assign n5520 = ~n964 ;
  assign n980 = n5520 & n979 ;
  assign n5521 = ~n949 ;
  assign n981 = n5521 & n980 ;
  assign n5522 = ~n297 ;
  assign n982 = n5522 & n981 ;
  assign n5523 = ~n253 ;
  assign n983 = n5523 & n982 ;
  assign n5524 = ~n256 ;
  assign n984 = n5524 & n983 ;
  assign n5525 = ~n552 ;
  assign n985 = n5525 & n984 ;
  assign n608 = n314 | n402 ;
  assign n609 = n473 | n608 ;
  assign n610 = n225 | n609 ;
  assign n611 = n345 | n610 ;
  assign n612 = n326 | n611 ;
  assign n613 = n151 | n612 ;
  assign n994 = n130 | n255 ;
  assign n995 = n365 | n994 ;
  assign n996 = n468 | n470 ;
  assign n997 = n995 | n996 ;
  assign n998 = n141 | n997 ;
  assign n999 = n324 | n998 ;
  assign n1000 = n445 | n999 ;
  assign n1001 = n312 | n1000 ;
  assign n1002 = n188 | n299 ;
  assign n1003 = n171 | n1002 ;
  assign n1004 = n189 | n1003 ;
  assign n1005 = n165 | n1004 ;
  assign n803 = n163 | n224 ;
  assign n1010 = n126 | n175 ;
  assign n1011 = n194 | n1010 ;
  assign n1012 = n448 | n1011 ;
  assign n1013 = n254 | n1012 ;
  assign n1014 = n1009 | n1013 ;
  assign n1015 = n952 | n1014 ;
  assign n1016 = n325 | n1015 ;
  assign n1017 = n173 | n1016 ;
  assign n1018 = n218 | n1017 ;
  assign n1019 = n169 | n1018 ;
  assign n1020 = n803 | n1019 ;
  assign n1021 = n221 | n1020 ;
  assign n1022 = n334 | n1021 ;
  assign n1023 = n172 | n1022 ;
  assign n1024 = n551 | n1023 ;
  assign n1025 = n348 | n1024 ;
  assign n1026 = n1005 | n1025 ;
  assign n1027 = n138 | n1026 ;
  assign n1028 = n1001 | n1027 ;
  assign n1029 = n993 | n1028 ;
  assign n1030 = n613 | n1029 ;
  assign n1031 = n296 | n1030 ;
  assign n1032 = n502 | n1031 ;
  assign n1033 = n364 | n1032 ;
  assign n5526 = ~n985 ;
  assign n1036 = n5526 & n1033 ;
  assign n5527 = ~n1036 ;
  assign n1037 = n802 & n5527 ;
  assign n1039 = n5473 & n5440 ;
  assign n1040 = x[7] & n1039 ;
  assign n1042 = x[7] | n1039 ;
  assign n5528 = ~n1040 ;
  assign n1043 = n5528 & n1042 ;
  assign n1044 = n441 & n1043 ;
  assign n5529 = ~n1037 ;
  assign n1045 = n5529 & n1044 ;
  assign n5530 = ~n1044 ;
  assign n1050 = n1037 & n5530 ;
  assign n1051 = n1045 | n1050 ;
  assign n5046 = x[8] & x[22] ;
  assign n5470 = x[8] & n5454 ;
  assign n847 = n5473 & n6771 ;
  assign n5531 = ~n5470 ;
  assign n849 = n5531 & n847 ;
  assign n1052 = n5046 | n849 ;
  assign n5532 = ~n1051 ;
  assign n1059 = n5532 & n1052 ;
  assign n1060 = n441 & n1059 ;
  assign n1061 = n1045 | n1060 ;
  assign n1063 = n931 & n1061 ;
  assign n4827 = x[14] & x[22] ;
  assign n57 = x[14] & n56 ;
  assign n5533 = ~n57 ;
  assign n521 = n5533 & n58 ;
  assign n522 = n5473 & n521 ;
  assign n523 = n4827 | n522 ;
  assign n577 = n114 | n194 ;
  assign n804 = n235 | n803 ;
  assign n805 = n476 | n804 ;
  assign n806 = n166 | n183 ;
  assign n807 = n344 | n806 ;
  assign n808 = n221 | n807 ;
  assign n646 = n124 | n325 ;
  assign n647 = n367 | n646 ;
  assign n811 = n131 | n175 ;
  assign n812 = n210 | n811 ;
  assign n813 = n810 | n812 ;
  assign n814 = n647 | n813 ;
  assign n815 = n808 | n814 ;
  assign n816 = n217 | n815 ;
  assign n817 = n347 | n816 ;
  assign n818 = n414 | n817 ;
  assign n819 = n130 | n818 ;
  assign n820 = n312 | n819 ;
  assign n821 = n101 | n820 ;
  assign n822 = n223 | n296 ;
  assign n823 = n120 | n172 ;
  assign n824 = n141 | n333 ;
  assign n323 = n5482 & n144 ;
  assign n614 = n150 | n429 ;
  assign n615 = n504 | n614 ;
  assign n616 = n613 | n615 ;
  assign n617 = n405 | n616 ;
  assign n618 = n186 | n617 ;
  assign n619 = n126 | n618 ;
  assign n620 = n215 | n619 ;
  assign n621 = n354 | n620 ;
  assign n622 = n323 | n621 ;
  assign n623 = n391 | n622 ;
  assign n624 = n348 | n623 ;
  assign n298 = n209 | n297 ;
  assign n825 = n457 | n588 ;
  assign n826 = n298 | n825 ;
  assign n827 = n146 | n826 ;
  assign n828 = n256 | n827 ;
  assign n829 = n365 | n828 ;
  assign n830 = n294 | n829 ;
  assign n831 = n204 | n830 ;
  assign n832 = n624 | n831 ;
  assign n833 = n824 | n832 ;
  assign n834 = n823 | n833 ;
  assign n835 = n822 | n834 ;
  assign n836 = n821 | n835 ;
  assign n837 = n805 | n836 ;
  assign n838 = n169 | n837 ;
  assign n839 = n577 | n838 ;
  assign n840 = n355 | n839 ;
  assign n841 = n752 | n840 ;
  assign n842 = n293 | n841 ;
  assign n5534 = ~n842 ;
  assign n843 = n802 & n5534 ;
  assign n5535 = ~n802 ;
  assign n889 = n5535 & n842 ;
  assign n890 = n843 | n889 ;
  assign n349 = n190 | n224 ;
  assign n350 = n348 | n349 ;
  assign n351 = n215 | n350 ;
  assign n352 = n214 | n351 ;
  assign n554 = n236 | n553 ;
  assign n555 = n206 | n554 ;
  assign n556 = n219 | n555 ;
  assign n557 = n364 | n556 ;
  assign n558 = n223 | n414 ;
  assign n559 = n293 | n558 ;
  assign n562 = n225 | n391 ;
  assign n563 = n124 | n562 ;
  assign n564 = n561 | n563 ;
  assign n565 = n559 | n564 ;
  assign n566 = n557 | n565 ;
  assign n567 = n182 | n566 ;
  assign n568 = n126 | n567 ;
  assign n569 = n345 | n568 ;
  assign n570 = n552 | n569 ;
  assign n573 = n334 | n572 ;
  assign n574 = n357 | n573 ;
  assign n575 = n210 | n574 ;
  assign n576 = n469 | n575 ;
  assign n578 = n110 | n577 ;
  assign n579 = n502 | n578 ;
  assign n580 = n468 | n579 ;
  assign n185 = n103 | n184 ;
  assign n581 = n170 & n185 ;
  assign n582 = n326 | n581 ;
  assign n583 = n448 | n582 ;
  assign n584 = n295 | n344 ;
  assign n585 = n353 | n584 ;
  assign n586 = n162 | n226 ;
  assign n587 = n356 | n586 ;
  assign n589 = n183 | n588 ;
  assign n590 = n587 | n589 ;
  assign n591 = n585 | n590 ;
  assign n592 = n583 | n591 ;
  assign n593 = n580 | n592 ;
  assign n594 = n576 | n593 ;
  assign n595 = n570 | n594 ;
  assign n596 = n352 | n595 ;
  assign n597 = n551 | n596 ;
  assign n844 = n802 | n842 ;
  assign n5536 = ~n597 ;
  assign n892 = n5536 & n844 ;
  assign n5537 = ~n892 ;
  assign n1064 = n890 & n5537 ;
  assign n1065 = n523 & n1064 ;
  assign n524 = n5473 & n55 ;
  assign n525 = x[13] & n524 ;
  assign n527 = x[13] | n524 ;
  assign n5538 = ~n525 ;
  assign n528 = n5538 & n527 ;
  assign n845 = n802 & n842 ;
  assign n5539 = ~n845 ;
  assign n846 = n597 & n5539 ;
  assign n891 = n846 | n890 ;
  assign n5540 = ~n528 ;
  assign n1075 = n5540 & n891 ;
  assign n893 = n890 | n892 ;
  assign n1085 = n528 & n893 ;
  assign n1086 = n1075 | n1085 ;
  assign n5541 = ~n846 ;
  assign n895 = n5541 & n890 ;
  assign n5542 = ~n523 ;
  assign n1087 = n5542 & n895 ;
  assign n5543 = ~n1087 ;
  assign n1088 = n1086 & n5543 ;
  assign n5544 = ~n1065 ;
  assign n1089 = n5544 & n1088 ;
  assign n4902 = x[12] & x[22] ;
  assign n54 = x[12] & n53 ;
  assign n5545 = ~n54 ;
  assign n526 = n5545 & n524 ;
  assign n677 = n4902 | n526 ;
  assign n359 = n357 | n358 ;
  assign n598 = n5482 & n113 ;
  assign n606 = n220 | n334 ;
  assign n607 = n110 | n606 ;
  assign n341 = n339 | n340 ;
  assign n625 = n206 | n212 ;
  assign n626 = n134 | n625 ;
  assign n627 = n166 | n626 ;
  assign n628 = n624 | n627 ;
  assign n629 = n341 | n628 ;
  assign n630 = n607 | n629 ;
  assign n631 = n605 | n630 ;
  assign n632 = n189 | n631 ;
  assign n633 = n445 | n632 ;
  assign n634 = n598 | n633 ;
  assign n635 = n209 | n634 ;
  assign n638 = n636 | n637 ;
  assign n639 = n194 | n638 ;
  assign n640 = n172 | n639 ;
  assign n641 = n297 | n640 ;
  assign n642 = n299 | n641 ;
  assign n643 = n211 | n471 ;
  assign n645 = n476 | n644 ;
  assign n648 = n254 | n647 ;
  assign n649 = n141 | n648 ;
  assign n650 = n219 | n649 ;
  assign n651 = n470 | n650 ;
  assign n652 = n129 | n651 ;
  assign n653 = n217 | n652 ;
  assign n654 = n457 | n653 ;
  assign n655 = n176 | n654 ;
  assign n656 = n645 | n655 ;
  assign n657 = n643 | n656 ;
  assign n658 = n642 | n657 ;
  assign n659 = n635 | n658 ;
  assign n660 = n359 | n659 ;
  assign n661 = n551 | n660 ;
  assign n662 = n364 | n661 ;
  assign n5546 = ~n662 ;
  assign n663 = n597 & n5546 ;
  assign n706 = n5536 & n662 ;
  assign n707 = n663 | n706 ;
  assign n664 = n597 | n662 ;
  assign n715 = n5507 & n664 ;
  assign n5547 = ~n715 ;
  assign n868 = n707 & n5547 ;
  assign n871 = n677 & n868 ;
  assign n665 = n597 & n662 ;
  assign n5548 = ~n665 ;
  assign n666 = n493 & n5548 ;
  assign n708 = n666 | n707 ;
  assign n712 = n5514 & n708 ;
  assign n716 = n707 | n715 ;
  assign n1090 = n672 & n716 ;
  assign n1091 = n712 | n1090 ;
  assign n5549 = ~n666 ;
  assign n717 = n5549 & n707 ;
  assign n5550 = ~n677 ;
  assign n1092 = n5550 & n717 ;
  assign n5551 = ~n1092 ;
  assign n1093 = n1091 & n5551 ;
  assign n5552 = ~n871 ;
  assign n1094 = n5552 & n1093 ;
  assign n1095 = n1089 & n1094 ;
  assign n862 = n685 & n859 ;
  assign n848 = x[9] & n847 ;
  assign n850 = x[9] | n847 ;
  assign n5553 = ~n848 ;
  assign n851 = n5553 & n850 ;
  assign n5554 = ~n851 ;
  assign n855 = n694 & n5554 ;
  assign n1096 = n543 & n851 ;
  assign n1097 = n855 | n1096 ;
  assign n1098 = n692 & n5512 ;
  assign n5555 = ~n1098 ;
  assign n1099 = n1097 & n5555 ;
  assign n5556 = ~n862 ;
  assign n1100 = n5556 & n1099 ;
  assign n1101 = n1089 | n1094 ;
  assign n5557 = ~n1095 ;
  assign n1102 = n5557 & n1101 ;
  assign n1104 = n1100 & n1102 ;
  assign n1105 = n1095 | n1104 ;
  assign n5558 = ~n1061 ;
  assign n1062 = n931 & n5558 ;
  assign n5559 = ~n931 ;
  assign n1106 = n5559 & n1061 ;
  assign n1107 = n1062 | n1106 ;
  assign n1109 = n1105 & n1107 ;
  assign n1110 = n1063 | n1109 ;
  assign n852 = n441 & n851 ;
  assign n853 = n5541 & n852 ;
  assign n5560 = ~n852 ;
  assign n857 = n846 & n5560 ;
  assign n858 = n853 | n857 ;
  assign n860 = n441 & n859 ;
  assign n5561 = ~n858 ;
  assign n861 = n5561 & n860 ;
  assign n5562 = ~n860 ;
  assign n1111 = n858 & n5562 ;
  assign n1112 = n861 | n1111 ;
  assign n5563 = ~n1112 ;
  assign n1114 = n1110 & n5563 ;
  assign n1113 = n1110 | n1112 ;
  assign n1115 = n1110 & n1112 ;
  assign n5564 = ~n1115 ;
  assign n1116 = n1113 & n5564 ;
  assign n5565 = ~n893 ;
  assign n894 = n523 & n5565 ;
  assign n896 = n523 | n846 ;
  assign n5566 = ~n895 ;
  assign n897 = n5566 & n896 ;
  assign n5567 = ~n894 ;
  assign n898 = n5567 & n897 ;
  assign n900 = n5560 & n898 ;
  assign n870 = n528 & n868 ;
  assign n711 = n5550 & n708 ;
  assign n901 = n677 & n716 ;
  assign n902 = n711 | n901 ;
  assign n903 = n5540 & n717 ;
  assign n5568 = ~n903 ;
  assign n904 = n902 & n5568 ;
  assign n5569 = ~n870 ;
  assign n905 = n5569 & n904 ;
  assign n899 = n852 & n898 ;
  assign n906 = n852 | n898 ;
  assign n5570 = ~n899 ;
  assign n907 = n5570 & n906 ;
  assign n5571 = ~n907 ;
  assign n908 = n905 & n5571 ;
  assign n909 = n900 | n908 ;
  assign n869 = n523 & n868 ;
  assign n709 = n5540 & n708 ;
  assign n878 = n528 & n716 ;
  assign n879 = n709 | n878 ;
  assign n880 = n5542 & n717 ;
  assign n5572 = ~n880 ;
  assign n881 = n879 & n5572 ;
  assign n5573 = ~n869 ;
  assign n882 = n5573 & n881 ;
  assign n689 = n677 & n685 ;
  assign n697 = n5514 & n694 ;
  assign n883 = n543 & n672 ;
  assign n884 = n697 | n883 ;
  assign n885 = n5550 & n692 ;
  assign n5574 = ~n885 ;
  assign n886 = n884 & n5574 ;
  assign n5575 = ~n689 ;
  assign n887 = n5575 & n886 ;
  assign n888 = n882 & n887 ;
  assign n910 = n882 | n887 ;
  assign n5576 = ~n888 ;
  assign n911 = n5576 & n910 ;
  assign n912 = n909 & n911 ;
  assign n1117 = n909 | n911 ;
  assign n5577 = ~n912 ;
  assign n1118 = n5577 & n1117 ;
  assign n5578 = ~n1116 ;
  assign n1119 = n5578 & n1118 ;
  assign n1120 = n1114 | n1119 ;
  assign n867 = n853 | n861 ;
  assign n913 = n888 | n912 ;
  assign n5579 = ~n913 ;
  assign n914 = n867 & n5579 ;
  assign n5580 = ~n867 ;
  assign n916 = n5580 & n913 ;
  assign n917 = n914 | n916 ;
  assign n688 = n528 & n685 ;
  assign n696 = n5550 & n694 ;
  assign n723 = n543 & n677 ;
  assign n724 = n696 | n723 ;
  assign n725 = n5540 & n692 ;
  assign n5581 = ~n725 ;
  assign n726 = n724 & n5581 ;
  assign n5582 = ~n688 ;
  assign n727 = n5582 & n726 ;
  assign n673 = n441 & n672 ;
  assign n667 = n523 | n666 ;
  assign n5583 = ~n717 ;
  assign n718 = n667 & n5583 ;
  assign n5584 = ~n716 ;
  assign n719 = n523 & n5584 ;
  assign n5585 = ~n719 ;
  assign n720 = n718 & n5585 ;
  assign n5586 = ~n720 ;
  assign n721 = n673 & n5586 ;
  assign n5587 = ~n673 ;
  assign n722 = n5587 & n720 ;
  assign n728 = n721 | n722 ;
  assign n5588 = ~n728 ;
  assign n729 = n727 & n5588 ;
  assign n5589 = ~n727 ;
  assign n918 = n5589 & n728 ;
  assign n919 = n729 | n918 ;
  assign n920 = n917 | n919 ;
  assign n1121 = n917 & n919 ;
  assign n5590 = ~n1121 ;
  assign n1122 = n920 & n5590 ;
  assign n5591 = ~n1122 ;
  assign n1124 = n1120 & n5591 ;
  assign n5592 = ~n1120 ;
  assign n1123 = n5592 & n1122 ;
  assign n1125 = n1123 | n1124 ;
  assign n872 = n672 & n868 ;
  assign n864 = n708 & n5512 ;
  assign n1126 = n716 & n859 ;
  assign n1127 = n864 | n1126 ;
  assign n1128 = n5514 & n717 ;
  assign n5593 = ~n1128 ;
  assign n1129 = n1127 & n5593 ;
  assign n5594 = ~n872 ;
  assign n1130 = n5594 & n1129 ;
  assign n854 = n685 & n851 ;
  assign n5595 = ~n1052 ;
  assign n1055 = n694 & n5595 ;
  assign n1131 = n543 & n1052 ;
  assign n1132 = n1055 | n1131 ;
  assign n1133 = n692 & n5554 ;
  assign n5596 = ~n1133 ;
  assign n1134 = n1132 & n5596 ;
  assign n5597 = ~n854 ;
  assign n1135 = n5597 & n1134 ;
  assign n1136 = n1130 & n1135 ;
  assign n301 = n176 | n300 ;
  assign n302 = n298 | n301 ;
  assign n303 = n134 | n302 ;
  assign n304 = n296 | n303 ;
  assign n305 = n189 | n304 ;
  assign n306 = n295 | n305 ;
  assign n307 = n294 | n306 ;
  assign n308 = n293 | n307 ;
  assign n1152 = n114 | n392 ;
  assign n1153 = n233 | n1152 ;
  assign n1154 = n447 | n1153 ;
  assign n1155 = n222 | n1154 ;
  assign n1156 = n459 | n467 ;
  assign n1157 = n173 | n1156 ;
  assign n1158 = n212 | n1157 ;
  assign n1159 = n216 | n1158 ;
  assign n1160 = n503 | n1159 ;
  assign n1161 = n355 | n1160 ;
  assign n1162 = n342 | n1161 ;
  assign n1163 = n221 | n598 ;
  assign n1164 = n137 | n333 ;
  assign n1165 = n1163 | n1164 ;
  assign n1166 = n608 | n1165 ;
  assign n1167 = n557 | n1166 ;
  assign n5598 = ~n1167 ;
  assign n1168 = n322 & n5598 ;
  assign n5599 = ~n1162 ;
  assign n1169 = n5599 & n1168 ;
  assign n5600 = ~n1155 ;
  assign n1170 = n5600 & n1169 ;
  assign n5601 = ~n308 ;
  assign n1171 = n5601 & n1170 ;
  assign n5602 = ~n1151 ;
  assign n1172 = n5602 & n1171 ;
  assign n5603 = ~n186 ;
  assign n1173 = n5603 & n1172 ;
  assign n5604 = ~n130 ;
  assign n1174 = n5604 & n1173 ;
  assign n5605 = ~n204 ;
  assign n1175 = n5605 & n1174 ;
  assign n5606 = ~n163 ;
  assign n1176 = n5606 & n1175 ;
  assign n5607 = ~n551 ;
  assign n1177 = n5607 & n1176 ;
  assign n1225 = n985 & n1177 ;
  assign n1179 = n458 | n1163 ;
  assign n1180 = n823 | n1179 ;
  assign n1181 = n218 | n1180 ;
  assign n1182 = n391 | n1181 ;
  assign n1183 = n645 | n974 ;
  assign n1184 = n311 | n1183 ;
  assign n1185 = n1155 | n1184 ;
  assign n1186 = n1182 | n1185 ;
  assign n1187 = n126 | n1186 ;
  assign n1188 = n194 | n1187 ;
  assign n1189 = n147 | n1188 ;
  assign n1190 = n211 | n1189 ;
  assign n1191 = n166 | n1190 ;
  assign n1192 = n312 | n1191 ;
  assign n1193 = n323 | n1192 ;
  assign n1194 = n636 | n937 ;
  assign n1195 = n192 | n1194 ;
  assign n1196 = n212 | n1195 ;
  assign n1197 = n345 | n1196 ;
  assign n1198 = n296 | n1197 ;
  assign n1199 = n551 | n1198 ;
  assign n1200 = n752 | n1199 ;
  assign n1201 = n559 | n995 ;
  assign n5608 = ~n1201 ;
  assign n1202 = n321 & n5608 ;
  assign n5609 = ~n1200 ;
  assign n1203 = n5609 & n1202 ;
  assign n5610 = ~n474 ;
  assign n1204 = n5610 & n1203 ;
  assign n5611 = ~n164 ;
  assign n1205 = n5611 & n1204 ;
  assign n5612 = ~n333 ;
  assign n1206 = n5612 & n1205 ;
  assign n1207 = n5524 & n1206 ;
  assign n5613 = ~n342 ;
  assign n1208 = n5613 & n1207 ;
  assign n5614 = ~n151 ;
  assign n1209 = n5614 & n1208 ;
  assign n5615 = ~n213 ;
  assign n1210 = n5615 & n1209 ;
  assign n360 = n356 | n359 ;
  assign n361 = n355 | n360 ;
  assign n362 = n354 | n361 ;
  assign n363 = n353 | n362 ;
  assign n1211 = n206 | n405 ;
  assign n1212 = n139 | n1211 ;
  assign n1213 = n108 | n1212 ;
  assign n1214 = n776 | n1213 ;
  assign n1215 = n450 | n1214 ;
  assign n1216 = n504 | n1215 ;
  assign n1217 = n363 | n1216 ;
  assign n1218 = n138 | n1217 ;
  assign n5616 = ~n1218 ;
  assign n1219 = n1210 & n5616 ;
  assign n5617 = ~n1193 ;
  assign n1220 = n5617 & n1219 ;
  assign n5618 = ~n149 ;
  assign n1221 = n5618 & n1220 ;
  assign n5619 = ~n217 ;
  assign n1222 = n5619 & n1221 ;
  assign n5620 = ~n332 ;
  assign n1223 = n5620 & n1222 ;
  assign n1226 = n1177 | n1223 ;
  assign n1227 = n5526 & n1226 ;
  assign n5621 = ~n1177 ;
  assign n1228 = n5621 & n1227 ;
  assign n5112 = x[6] & x[22] ;
  assign n5424 = x[6] & n5401 ;
  assign n5622 = ~n5424 ;
  assign n1041 = n5622 & n1039 ;
  assign n1229 = n5112 | n1041 ;
  assign n1230 = n441 & n1229 ;
  assign n5623 = ~n1225 ;
  assign n1239 = n5623 & n1230 ;
  assign n5624 = ~n1228 ;
  assign n1240 = n5624 & n1239 ;
  assign n1242 = n1225 | n1240 ;
  assign n1244 = n1130 | n1135 ;
  assign n5625 = ~n1136 ;
  assign n1245 = n5625 & n1244 ;
  assign n1247 = n1242 & n1245 ;
  assign n1248 = n1136 | n1247 ;
  assign n1038 = n523 | n1037 ;
  assign n1034 = n985 | n1033 ;
  assign n1249 = n985 & n1033 ;
  assign n5626 = ~n1249 ;
  assign n1250 = n1034 & n5626 ;
  assign n1265 = n1037 | n1250 ;
  assign n1274 = n1038 & n1265 ;
  assign n5627 = ~n1033 ;
  assign n1035 = n985 & n5627 ;
  assign n1263 = n802 | n1035 ;
  assign n1264 = n1250 & n1263 ;
  assign n1275 = n523 & n1264 ;
  assign n5628 = ~n1275 ;
  assign n1276 = n1274 & n5628 ;
  assign n1278 = n5530 & n1276 ;
  assign n1066 = n528 & n1064 ;
  assign n1077 = n5550 & n891 ;
  assign n1279 = n677 & n893 ;
  assign n1280 = n1077 | n1279 ;
  assign n1281 = n5540 & n895 ;
  assign n5629 = ~n1281 ;
  assign n1282 = n1280 & n5629 ;
  assign n5630 = ~n1066 ;
  assign n1283 = n5630 & n1282 ;
  assign n5631 = ~n1276 ;
  assign n1277 = n1044 & n5631 ;
  assign n1284 = n1277 | n1278 ;
  assign n5632 = ~n1284 ;
  assign n1285 = n1283 & n5632 ;
  assign n1286 = n1278 | n1285 ;
  assign n1288 = n1248 & n1286 ;
  assign n1287 = n1248 | n1286 ;
  assign n5633 = ~n1288 ;
  assign n1289 = n1287 & n5633 ;
  assign n5634 = ~n1059 ;
  assign n1290 = n441 & n5634 ;
  assign n1291 = n1052 & n1290 ;
  assign n1292 = n1051 | n1060 ;
  assign n5635 = ~n1291 ;
  assign n1293 = n5635 & n1292 ;
  assign n5636 = ~n1293 ;
  assign n1295 = n1289 & n5636 ;
  assign n1296 = n1288 | n1295 ;
  assign n5637 = ~n905 ;
  assign n1297 = n5637 & n907 ;
  assign n1298 = n908 | n1297 ;
  assign n5638 = ~n1298 ;
  assign n1300 = n1296 & n5638 ;
  assign n1108 = n1105 | n1107 ;
  assign n5639 = ~n1109 ;
  assign n1301 = n1108 & n5639 ;
  assign n1299 = n1296 | n1298 ;
  assign n1302 = n1296 & n1298 ;
  assign n5640 = ~n1302 ;
  assign n1303 = n1299 & n5640 ;
  assign n5641 = ~n1303 ;
  assign n1304 = n1301 & n5641 ;
  assign n1306 = n1300 | n1304 ;
  assign n5642 = ~n1118 ;
  assign n1307 = n1116 & n5642 ;
  assign n1308 = n1119 | n1307 ;
  assign n5643 = ~n1308 ;
  assign n1310 = n1306 & n5643 ;
  assign n1305 = n1301 | n1303 ;
  assign n1311 = n1301 & n1303 ;
  assign n5644 = ~n1311 ;
  assign n1312 = n1305 & n5644 ;
  assign n873 = n859 & n868 ;
  assign n856 = n708 & n5554 ;
  assign n1313 = n716 & n851 ;
  assign n1314 = n856 | n1313 ;
  assign n1315 = n717 & n5512 ;
  assign n5645 = ~n1315 ;
  assign n1316 = n1314 & n5645 ;
  assign n5646 = ~n873 ;
  assign n1317 = n5646 & n1316 ;
  assign n1053 = n685 & n1052 ;
  assign n5647 = ~n1043 ;
  assign n1047 = n694 & n5647 ;
  assign n1318 = n543 & n1043 ;
  assign n1319 = n1047 | n1318 ;
  assign n1320 = n692 & n5595 ;
  assign n5648 = ~n1320 ;
  assign n1321 = n1319 & n5648 ;
  assign n5649 = ~n1053 ;
  assign n1322 = n5649 & n1321 ;
  assign n1323 = n1317 & n1322 ;
  assign n1266 = n523 | n1265 ;
  assign n1251 = n5529 & n1250 ;
  assign n1255 = n5540 & n1251 ;
  assign n1328 = n528 & n1264 ;
  assign n1329 = n1255 | n1328 ;
  assign n5650 = ~n1329 ;
  assign n1330 = n1266 & n5650 ;
  assign n5651 = ~n1250 ;
  assign n1324 = n5651 & n1263 ;
  assign n1331 = n523 & n1324 ;
  assign n5652 = ~n1331 ;
  assign n1332 = n1330 & n5652 ;
  assign n1333 = n1317 | n1322 ;
  assign n5653 = ~n1323 ;
  assign n1334 = n5653 & n1333 ;
  assign n1336 = n1332 & n1334 ;
  assign n1337 = n1323 | n1336 ;
  assign n5654 = ~n1283 ;
  assign n1338 = n5654 & n1284 ;
  assign n1339 = n1285 | n1338 ;
  assign n5655 = ~n1339 ;
  assign n1341 = n1337 & n5655 ;
  assign n1340 = n1337 | n1339 ;
  assign n1342 = n1337 & n1339 ;
  assign n5656 = ~n1342 ;
  assign n1343 = n1340 & n5656 ;
  assign n5657 = ~n1242 ;
  assign n1246 = n5657 & n1245 ;
  assign n5658 = ~n1245 ;
  assign n1344 = n1242 & n5658 ;
  assign n1345 = n1246 | n1344 ;
  assign n5659 = ~n1343 ;
  assign n1347 = n5659 & n1345 ;
  assign n1348 = n1341 | n1347 ;
  assign n5660 = ~n1102 ;
  assign n1103 = n1100 & n5660 ;
  assign n5661 = ~n1100 ;
  assign n1349 = n5661 & n1102 ;
  assign n1350 = n1103 | n1349 ;
  assign n1352 = n1348 & n1350 ;
  assign n1351 = n1348 | n1350 ;
  assign n5662 = ~n1352 ;
  assign n1353 = n1351 & n5662 ;
  assign n5663 = ~n1289 ;
  assign n1294 = n5663 & n1293 ;
  assign n1354 = n1294 | n1295 ;
  assign n5664 = ~n1354 ;
  assign n1355 = n1353 & n5664 ;
  assign n1357 = n1352 | n1355 ;
  assign n5665 = ~n1312 ;
  assign n1359 = n5665 & n1357 ;
  assign n5666 = ~n1357 ;
  assign n1358 = n1312 & n5666 ;
  assign n1360 = n1358 | n1359 ;
  assign n1067 = n677 & n1064 ;
  assign n1079 = n5514 & n891 ;
  assign n1361 = n672 & n893 ;
  assign n1362 = n1079 | n1361 ;
  assign n1363 = n5550 & n895 ;
  assign n5667 = ~n1363 ;
  assign n1364 = n1362 & n5667 ;
  assign n5668 = ~n1067 ;
  assign n1365 = n5668 & n1364 ;
  assign n5669 = ~n1240 ;
  assign n1241 = n1230 & n5669 ;
  assign n1243 = n1228 | n1242 ;
  assign n5670 = ~n1241 ;
  assign n1366 = n5670 & n1243 ;
  assign n5671 = ~n1366 ;
  assign n1368 = n1365 & n5671 ;
  assign n443 = n274 & n441 ;
  assign n1370 = n443 & n5621 ;
  assign n5672 = ~n443 ;
  assign n1369 = n5672 & n1177 ;
  assign n1224 = n1177 & n1223 ;
  assign n5673 = ~n1224 ;
  assign n1372 = n5673 & n1226 ;
  assign n5674 = ~n1372 ;
  assign n1386 = n523 & n5674 ;
  assign n1387 = n1227 | n1386 ;
  assign n1384 = n985 & n5673 ;
  assign n1385 = n1372 | n1384 ;
  assign n5675 = ~n1385 ;
  assign n1388 = n523 & n5675 ;
  assign n5676 = ~n1388 ;
  assign n1389 = n1387 & n5676 ;
  assign n5677 = ~n1369 ;
  assign n1390 = n5677 & n1389 ;
  assign n1391 = n1370 | n1390 ;
  assign n1367 = n1365 & n1366 ;
  assign n1392 = n1365 | n1366 ;
  assign n5678 = ~n1367 ;
  assign n1393 = n5678 & n1392 ;
  assign n5679 = ~n1393 ;
  assign n1394 = n1391 & n5679 ;
  assign n1395 = n1368 | n1394 ;
  assign n1268 = n528 | n1265 ;
  assign n1257 = n5550 & n1251 ;
  assign n1396 = n677 & n1264 ;
  assign n1397 = n1257 | n1396 ;
  assign n5680 = ~n1397 ;
  assign n1398 = n1268 & n5680 ;
  assign n1399 = n528 & n1324 ;
  assign n5681 = ~n1399 ;
  assign n1400 = n1398 & n5681 ;
  assign n1071 = n672 & n1064 ;
  assign n1080 = n5512 & n891 ;
  assign n1401 = n859 & n893 ;
  assign n1402 = n1080 | n1401 ;
  assign n1403 = n5514 & n895 ;
  assign n5682 = ~n1403 ;
  assign n1404 = n1402 & n5682 ;
  assign n5683 = ~n1071 ;
  assign n1405 = n5683 & n1404 ;
  assign n1407 = n1400 & n1405 ;
  assign n874 = n851 & n868 ;
  assign n1056 = n708 & n5595 ;
  assign n1408 = n716 & n1052 ;
  assign n1409 = n1056 | n1408 ;
  assign n1410 = n717 & n5554 ;
  assign n5684 = ~n1410 ;
  assign n1411 = n1409 & n5684 ;
  assign n5685 = ~n874 ;
  assign n1412 = n5685 & n1411 ;
  assign n5686 = ~n1400 ;
  assign n1406 = n5686 & n1405 ;
  assign n5687 = ~n1405 ;
  assign n1413 = n1400 & n5687 ;
  assign n1414 = n1406 | n1413 ;
  assign n1416 = n1412 & n1414 ;
  assign n1417 = n1407 | n1416 ;
  assign n1335 = n1332 | n1334 ;
  assign n5688 = ~n1336 ;
  assign n1418 = n1335 & n5688 ;
  assign n1419 = n1417 & n1418 ;
  assign n1048 = n692 & n5647 ;
  assign n1234 = n694 | n1229 ;
  assign n5689 = ~n543 ;
  assign n1420 = n5689 & n1229 ;
  assign n5690 = ~n1420 ;
  assign n1421 = n1234 & n5690 ;
  assign n5691 = ~n1048 ;
  assign n1422 = n5691 & n1421 ;
  assign n1423 = n685 & n1043 ;
  assign n5692 = ~n1423 ;
  assign n1424 = n1422 & n5692 ;
  assign n442 = n275 & n441 ;
  assign n1426 = n442 & n5621 ;
  assign n5693 = ~n442 ;
  assign n1425 = n5693 & n1177 ;
  assign n5694 = ~n1384 ;
  assign n1428 = n1372 & n5694 ;
  assign n1433 = n523 & n1428 ;
  assign n1373 = n1227 | n1372 ;
  assign n1374 = n5540 & n1373 ;
  assign n1441 = n528 & n1385 ;
  assign n1442 = n1374 | n1441 ;
  assign n5695 = ~n1227 ;
  assign n1434 = n5695 & n1372 ;
  assign n1443 = n5542 & n1434 ;
  assign n5696 = ~n1443 ;
  assign n1444 = n1442 & n5696 ;
  assign n5697 = ~n1433 ;
  assign n1445 = n5697 & n1444 ;
  assign n5698 = ~n1425 ;
  assign n1446 = n5698 & n1445 ;
  assign n1447 = n1426 | n1446 ;
  assign n1450 = n1424 & n1447 ;
  assign n1448 = n1424 | n1447 ;
  assign n5699 = ~n1450 ;
  assign n1451 = n1448 & n5699 ;
  assign n1068 = n859 & n1064 ;
  assign n1081 = n5554 & n891 ;
  assign n1452 = n851 & n893 ;
  assign n1453 = n1081 | n1452 ;
  assign n1454 = n5512 & n895 ;
  assign n5700 = ~n1454 ;
  assign n1455 = n1453 & n5700 ;
  assign n5701 = ~n1068 ;
  assign n1456 = n5701 & n1455 ;
  assign n1325 = n677 & n1324 ;
  assign n1252 = n672 | n1251 ;
  assign n5702 = ~n1264 ;
  assign n1457 = n672 & n5702 ;
  assign n5703 = ~n1457 ;
  assign n1458 = n1252 & n5703 ;
  assign n1459 = n677 | n1265 ;
  assign n5704 = ~n1458 ;
  assign n1460 = n5704 & n1459 ;
  assign n5705 = ~n1325 ;
  assign n1461 = n5705 & n1460 ;
  assign n1462 = n1456 & n1461 ;
  assign n1054 = n868 & n1052 ;
  assign n1049 = n708 & n5647 ;
  assign n1463 = n716 & n1043 ;
  assign n1464 = n1049 | n1463 ;
  assign n1465 = n717 & n5595 ;
  assign n5706 = ~n1465 ;
  assign n1466 = n1464 & n5706 ;
  assign n5707 = ~n1054 ;
  assign n1467 = n5707 & n1466 ;
  assign n1468 = n1456 | n1461 ;
  assign n5708 = ~n1462 ;
  assign n1469 = n5708 & n1468 ;
  assign n1471 = n1467 & n1469 ;
  assign n1472 = n1462 | n1471 ;
  assign n1474 = n1451 & n1472 ;
  assign n1475 = n1450 | n1474 ;
  assign n1476 = n1417 | n1418 ;
  assign n5709 = ~n1419 ;
  assign n1477 = n5709 & n1476 ;
  assign n1478 = n1475 & n1477 ;
  assign n1479 = n1419 | n1478 ;
  assign n1481 = n1395 & n1479 ;
  assign n1480 = n1395 | n1479 ;
  assign n5710 = ~n1481 ;
  assign n1482 = n1480 & n5710 ;
  assign n1346 = n1343 & n1345 ;
  assign n1483 = n1343 | n1345 ;
  assign n5711 = ~n1346 ;
  assign n1484 = n5711 & n1483 ;
  assign n5712 = ~n1484 ;
  assign n1486 = n1482 & n5712 ;
  assign n1487 = n1481 | n1486 ;
  assign n1356 = n1353 & n1354 ;
  assign n1488 = n1353 | n1354 ;
  assign n5713 = ~n1356 ;
  assign n1489 = n5713 & n1488 ;
  assign n5714 = ~n1489 ;
  assign n1491 = n1487 & n5714 ;
  assign n5715 = ~n1482 ;
  assign n1485 = n5715 & n1484 ;
  assign n1492 = n1485 | n1486 ;
  assign n1493 = n1369 | n1391 ;
  assign n1371 = n1369 | n1370 ;
  assign n1494 = n1371 & n1389 ;
  assign n5716 = ~n1494 ;
  assign n1495 = n1493 & n5716 ;
  assign n5717 = ~n1414 ;
  assign n1415 = n1412 & n5717 ;
  assign n5718 = ~n1412 ;
  assign n1496 = n5718 & n1414 ;
  assign n1497 = n1415 | n1496 ;
  assign n5719 = ~n1495 ;
  assign n1499 = n5719 & n1497 ;
  assign n5720 = ~n1497 ;
  assign n1498 = n1495 & n5720 ;
  assign n1500 = n1498 | n1499 ;
  assign n1231 = n685 & n1229 ;
  assign n5721 = ~n274 ;
  assign n699 = n5721 & n694 ;
  assign n1501 = n274 & n543 ;
  assign n1502 = n699 | n1501 ;
  assign n5722 = ~n1229 ;
  assign n1503 = n692 & n5722 ;
  assign n5723 = ~n1503 ;
  assign n1504 = n1502 & n5723 ;
  assign n5724 = ~n1231 ;
  assign n1505 = n5724 & n1504 ;
  assign n1506 = n282 & n441 ;
  assign n1507 = n219 | n825 ;
  assign n1508 = n171 | n1507 ;
  assign n1509 = n297 | n1508 ;
  assign n1510 = n120 | n1509 ;
  assign n1511 = n210 | n1510 ;
  assign n1512 = n344 | n1511 ;
  assign n1513 = n551 | n1512 ;
  assign n1514 = n552 | n1513 ;
  assign n1515 = n218 | n347 ;
  assign n1516 = n312 | n1515 ;
  assign n1517 = n429 | n583 ;
  assign n1518 = n1516 | n1517 ;
  assign n1519 = n994 | n1518 ;
  assign n1520 = n643 | n1519 ;
  assign n1521 = n334 | n1520 ;
  assign n1522 = n212 | n1521 ;
  assign n1523 = n414 | n1522 ;
  assign n1524 = n232 | n1523 ;
  assign n1525 = n364 | n1524 ;
  assign n5725 = ~n357 ;
  assign n1526 = n321 & n5725 ;
  assign n5726 = ~n445 ;
  assign n1527 = n5726 & n1526 ;
  assign n5727 = ~n169 ;
  assign n1528 = n5727 & n1527 ;
  assign n5728 = ~n502 ;
  assign n1529 = n5728 & n1528 ;
  assign n5729 = ~n353 ;
  assign n1530 = n5729 & n1529 ;
  assign n5730 = ~n214 ;
  assign n1531 = n5730 & n1530 ;
  assign n5731 = ~n339 ;
  assign n1532 = n5731 & n1531 ;
  assign n1533 = n5614 & n1532 ;
  assign n5732 = ~n370 ;
  assign n1534 = n5732 & n1533 ;
  assign n5733 = ~n1525 ;
  assign n1535 = n5733 & n1534 ;
  assign n5734 = ~n418 ;
  assign n1536 = n5734 & n1535 ;
  assign n5735 = ~n1514 ;
  assign n1537 = n5735 & n1536 ;
  assign n5736 = ~n175 ;
  assign n1538 = n5736 & n1537 ;
  assign n5737 = ~n206 ;
  assign n1539 = n5737 & n1538 ;
  assign n5738 = ~n114 ;
  assign n1540 = n5738 & n1539 ;
  assign n5739 = ~n358 ;
  assign n1541 = n5739 & n1540 ;
  assign n1542 = n5524 & n1541 ;
  assign n5740 = ~n598 ;
  assign n1543 = n5740 & n1542 ;
  assign n5741 = ~n209 ;
  assign n1544 = n5741 & n1543 ;
  assign n1547 = n523 & n1544 ;
  assign n1548 = n1177 | n1547 ;
  assign n5742 = ~n1548 ;
  assign n1550 = n1506 & n5742 ;
  assign n1429 = n528 & n1428 ;
  assign n1376 = n5550 & n1373 ;
  assign n1551 = n677 & n1385 ;
  assign n1552 = n1376 | n1551 ;
  assign n1553 = n5540 & n1434 ;
  assign n5743 = ~n1553 ;
  assign n1554 = n1552 & n5743 ;
  assign n5744 = ~n1429 ;
  assign n1555 = n5744 & n1554 ;
  assign n1549 = n1506 & n1548 ;
  assign n1556 = n1506 | n1548 ;
  assign n5745 = ~n1549 ;
  assign n1557 = n5745 & n1556 ;
  assign n5746 = ~n1557 ;
  assign n1558 = n1555 & n5746 ;
  assign n1559 = n1550 | n1558 ;
  assign n1561 = n1505 & n1559 ;
  assign n5747 = ~n1559 ;
  assign n1560 = n1505 & n5747 ;
  assign n5748 = ~n1505 ;
  assign n1562 = n5748 & n1559 ;
  assign n1563 = n1560 | n1562 ;
  assign n1069 = n851 & n1064 ;
  assign n1078 = n891 & n5595 ;
  assign n1564 = n893 & n1052 ;
  assign n1565 = n1078 | n1564 ;
  assign n1566 = n5554 & n895 ;
  assign n5749 = ~n1566 ;
  assign n1567 = n1565 & n5749 ;
  assign n5750 = ~n1069 ;
  assign n1568 = n5750 & n1567 ;
  assign n1326 = n672 & n1324 ;
  assign n1253 = n859 | n1251 ;
  assign n1569 = n859 & n5702 ;
  assign n5751 = ~n1569 ;
  assign n1570 = n1253 & n5751 ;
  assign n1571 = n672 | n1265 ;
  assign n5752 = ~n1570 ;
  assign n1572 = n5752 & n1571 ;
  assign n5753 = ~n1326 ;
  assign n1573 = n5753 & n1572 ;
  assign n1574 = n1568 & n1573 ;
  assign n1046 = n868 & n1043 ;
  assign n1235 = n708 & n5722 ;
  assign n1575 = n716 & n1229 ;
  assign n1576 = n1235 | n1575 ;
  assign n1577 = n717 & n5647 ;
  assign n5754 = ~n1577 ;
  assign n1578 = n1576 & n5754 ;
  assign n5755 = ~n1046 ;
  assign n1579 = n5755 & n1578 ;
  assign n1580 = n1568 | n1573 ;
  assign n5756 = ~n1574 ;
  assign n1581 = n5756 & n1580 ;
  assign n1583 = n1579 & n1581 ;
  assign n1584 = n1574 | n1583 ;
  assign n1586 = n1563 & n1584 ;
  assign n1587 = n1561 | n1586 ;
  assign n5757 = ~n1500 ;
  assign n1589 = n5757 & n1587 ;
  assign n1590 = n1499 | n1589 ;
  assign n5758 = ~n1391 ;
  assign n1591 = n5758 & n1393 ;
  assign n1592 = n1394 | n1591 ;
  assign n5759 = ~n1592 ;
  assign n1593 = n1590 & n5759 ;
  assign n5760 = ~n1590 ;
  assign n1594 = n5760 & n1592 ;
  assign n1595 = n1593 | n1594 ;
  assign n1596 = n1475 | n1477 ;
  assign n5761 = ~n1478 ;
  assign n1597 = n5761 & n1596 ;
  assign n5762 = ~n1595 ;
  assign n1598 = n5762 & n1597 ;
  assign n1599 = n1593 | n1598 ;
  assign n5763 = ~n1492 ;
  assign n1601 = n5763 & n1599 ;
  assign n5764 = ~n1599 ;
  assign n1600 = n1492 & n5764 ;
  assign n1602 = n1600 | n1601 ;
  assign n1603 = n1177 | n1544 ;
  assign n5765 = ~n1603 ;
  assign n1604 = n523 & n5765 ;
  assign n5766 = ~n1544 ;
  assign n1545 = n1177 & n5766 ;
  assign n1613 = n5542 & n1545 ;
  assign n1612 = n528 | n1177 ;
  assign n1614 = n1544 & n1612 ;
  assign n1615 = n1613 | n1614 ;
  assign n1616 = n1604 | n1615 ;
  assign n691 = n282 & n685 ;
  assign n539 = n282 & n538 ;
  assign n1617 = n539 | n545 ;
  assign n5767 = ~n691 ;
  assign n1618 = n5767 & n1617 ;
  assign n1619 = n545 & n1618 ;
  assign n5768 = ~n1616 ;
  assign n1620 = n5768 & n1619 ;
  assign n690 = n274 & n685 ;
  assign n698 = n5498 & n694 ;
  assign n1621 = n275 & n543 ;
  assign n1622 = n698 | n1621 ;
  assign n1623 = n5721 & n692 ;
  assign n5769 = ~n1623 ;
  assign n1624 = n1622 & n5769 ;
  assign n5770 = ~n690 ;
  assign n1625 = n5770 & n1624 ;
  assign n1626 = n1620 & n1625 ;
  assign n1072 = n1052 & n1064 ;
  assign n1082 = n891 & n5647 ;
  assign n1627 = n893 & n1043 ;
  assign n1628 = n1082 | n1627 ;
  assign n1629 = n895 & n5595 ;
  assign n5771 = ~n1629 ;
  assign n1630 = n1628 & n5771 ;
  assign n5772 = ~n1072 ;
  assign n1631 = n5772 & n1630 ;
  assign n1232 = n868 & n1229 ;
  assign n713 = n5721 & n708 ;
  assign n1632 = n274 & n716 ;
  assign n1633 = n713 | n1632 ;
  assign n1634 = n717 & n5722 ;
  assign n5773 = ~n1634 ;
  assign n1635 = n1633 & n5773 ;
  assign n5774 = ~n1232 ;
  assign n1636 = n5774 & n1635 ;
  assign n1637 = n1631 & n1636 ;
  assign n1270 = n859 | n1265 ;
  assign n1258 = n5554 & n1251 ;
  assign n1638 = n851 & n1264 ;
  assign n1639 = n1258 | n1638 ;
  assign n5775 = ~n1639 ;
  assign n1640 = n1270 & n5775 ;
  assign n1641 = n859 & n1324 ;
  assign n5776 = ~n1641 ;
  assign n1642 = n1640 & n5776 ;
  assign n1643 = n1631 | n1636 ;
  assign n5777 = ~n1637 ;
  assign n1644 = n5777 & n1643 ;
  assign n1646 = n1642 & n1644 ;
  assign n1647 = n1637 | n1646 ;
  assign n1648 = n1620 | n1625 ;
  assign n5778 = ~n1626 ;
  assign n1649 = n5778 & n1648 ;
  assign n1651 = n1647 & n1649 ;
  assign n1652 = n1626 | n1651 ;
  assign n1449 = n1425 | n1447 ;
  assign n1427 = n1425 | n1426 ;
  assign n1653 = n1427 & n1445 ;
  assign n5779 = ~n1653 ;
  assign n1654 = n1449 & n5779 ;
  assign n5780 = ~n1654 ;
  assign n1661 = n1652 & n5780 ;
  assign n1655 = n1652 & n1654 ;
  assign n1656 = n1652 | n1654 ;
  assign n5781 = ~n1655 ;
  assign n1657 = n5781 & n1656 ;
  assign n5782 = ~n1469 ;
  assign n1470 = n1467 & n5782 ;
  assign n5783 = ~n1467 ;
  assign n1658 = n5783 & n1469 ;
  assign n1659 = n1470 | n1658 ;
  assign n5784 = ~n1657 ;
  assign n1662 = n5784 & n1659 ;
  assign n1663 = n1661 | n1662 ;
  assign n1473 = n1451 | n1472 ;
  assign n5785 = ~n1474 ;
  assign n1664 = n1473 & n5785 ;
  assign n1665 = n1663 & n1664 ;
  assign n5786 = ~n1587 ;
  assign n1588 = n1500 & n5786 ;
  assign n1666 = n1588 | n1589 ;
  assign n1667 = n1663 | n1664 ;
  assign n5787 = ~n1665 ;
  assign n1668 = n5787 & n1667 ;
  assign n5788 = ~n1666 ;
  assign n1670 = n5788 & n1668 ;
  assign n1671 = n1665 | n1670 ;
  assign n5789 = ~n1597 ;
  assign n1672 = n1595 & n5789 ;
  assign n1673 = n1598 | n1672 ;
  assign n5790 = ~n1673 ;
  assign n1675 = n1671 & n5790 ;
  assign n1435 = n5550 & n1434 ;
  assign n1379 = n672 | n1373 ;
  assign n1676 = n672 & n5675 ;
  assign n5791 = ~n1676 ;
  assign n1677 = n1379 & n5791 ;
  assign n5792 = ~n1435 ;
  assign n1678 = n5792 & n1677 ;
  assign n1679 = n677 & n1428 ;
  assign n5793 = ~n1679 ;
  assign n1680 = n1678 & n5793 ;
  assign n693 = n5498 & n692 ;
  assign n700 = n282 | n694 ;
  assign n1681 = n282 & n5689 ;
  assign n5794 = ~n1681 ;
  assign n1682 = n700 & n5794 ;
  assign n5795 = ~n693 ;
  assign n1683 = n5795 & n1682 ;
  assign n1684 = n275 & n685 ;
  assign n5796 = ~n1684 ;
  assign n1685 = n1683 & n5796 ;
  assign n1687 = n1680 & n1685 ;
  assign n1686 = n1680 | n1685 ;
  assign n5797 = ~n1619 ;
  assign n1688 = n1616 & n5797 ;
  assign n1689 = n1620 | n1688 ;
  assign n5798 = ~n1689 ;
  assign n1690 = n1686 & n5798 ;
  assign n1691 = n1687 | n1690 ;
  assign n5799 = ~n1555 ;
  assign n1693 = n5799 & n1557 ;
  assign n1694 = n1558 | n1693 ;
  assign n5800 = ~n1694 ;
  assign n1696 = n1691 & n5800 ;
  assign n1695 = n1691 | n1694 ;
  assign n1697 = n1691 & n1694 ;
  assign n5801 = ~n1697 ;
  assign n1698 = n1695 & n5801 ;
  assign n5802 = ~n1581 ;
  assign n1582 = n1579 & n5802 ;
  assign n5803 = ~n1579 ;
  assign n1699 = n5803 & n1581 ;
  assign n1700 = n1582 | n1699 ;
  assign n5804 = ~n1698 ;
  assign n1702 = n5804 & n1700 ;
  assign n1703 = n1696 | n1702 ;
  assign n5805 = ~n1584 ;
  assign n1585 = n1563 & n5805 ;
  assign n5806 = ~n1563 ;
  assign n1704 = n5806 & n1584 ;
  assign n1705 = n1585 | n1704 ;
  assign n1707 = n1703 & n1705 ;
  assign n5807 = ~n1703 ;
  assign n1706 = n5807 & n1705 ;
  assign n5808 = ~n1705 ;
  assign n1708 = n1703 & n5808 ;
  assign n1709 = n1706 | n1708 ;
  assign n5809 = ~n1659 ;
  assign n1660 = n1657 & n5809 ;
  assign n1710 = n1660 | n1662 ;
  assign n5810 = ~n1710 ;
  assign n1711 = n1709 & n5810 ;
  assign n1712 = n1707 | n1711 ;
  assign n1669 = n1666 & n1668 ;
  assign n1713 = n1666 | n1668 ;
  assign n5811 = ~n1669 ;
  assign n1714 = n5811 & n1713 ;
  assign n5812 = ~n1714 ;
  assign n1716 = n1712 & n5812 ;
  assign n1272 = n851 | n1265 ;
  assign n1259 = n5595 & n1251 ;
  assign n1728 = n1052 & n1264 ;
  assign n1729 = n1259 | n1728 ;
  assign n5813 = ~n1729 ;
  assign n1730 = n1272 & n5813 ;
  assign n1731 = n851 & n1324 ;
  assign n5814 = ~n1731 ;
  assign n1732 = n1730 & n5814 ;
  assign n1073 = n1043 & n1064 ;
  assign n1236 = n891 & n5722 ;
  assign n1733 = n893 & n1229 ;
  assign n1734 = n1236 | n1733 ;
  assign n1735 = n895 & n5647 ;
  assign n5815 = ~n1735 ;
  assign n1736 = n1734 & n5815 ;
  assign n5816 = ~n1073 ;
  assign n1737 = n5816 & n1736 ;
  assign n1742 = n1732 & n1737 ;
  assign n1605 = n677 & n5765 ;
  assign n1718 = n5550 & n1545 ;
  assign n1717 = n672 | n1177 ;
  assign n1719 = n1544 & n1717 ;
  assign n1720 = n1718 | n1719 ;
  assign n1721 = n1605 | n1720 ;
  assign n875 = n282 & n868 ;
  assign n1722 = n282 & n707 ;
  assign n1723 = n666 | n1722 ;
  assign n5817 = ~n875 ;
  assign n1724 = n5817 & n1723 ;
  assign n1725 = n666 & n1724 ;
  assign n5818 = ~n1721 ;
  assign n1727 = n5818 & n1725 ;
  assign n5819 = ~n1732 ;
  assign n1738 = n5819 & n1737 ;
  assign n5820 = ~n1737 ;
  assign n1739 = n1732 & n5820 ;
  assign n1740 = n1738 | n1739 ;
  assign n1743 = n1727 & n1740 ;
  assign n1744 = n1742 | n1743 ;
  assign n1606 = n528 & n5765 ;
  assign n1746 = n5540 & n1545 ;
  assign n1745 = n677 | n1177 ;
  assign n1747 = n1544 & n1745 ;
  assign n1748 = n1746 | n1747 ;
  assign n1749 = n1606 | n1748 ;
  assign n1430 = n672 & n1428 ;
  assign n1377 = n5512 & n1373 ;
  assign n1750 = n859 & n1385 ;
  assign n1751 = n1377 | n1750 ;
  assign n1752 = n5514 & n1434 ;
  assign n5821 = ~n1752 ;
  assign n1753 = n1751 & n5821 ;
  assign n5822 = ~n1430 ;
  assign n1754 = n5822 & n1753 ;
  assign n5823 = ~n1749 ;
  assign n1755 = n5823 & n1754 ;
  assign n876 = n274 & n868 ;
  assign n710 = n5498 & n708 ;
  assign n1756 = n275 & n716 ;
  assign n1757 = n710 | n1756 ;
  assign n1758 = n5721 & n717 ;
  assign n5824 = ~n1758 ;
  assign n1759 = n1757 & n5824 ;
  assign n5825 = ~n876 ;
  assign n1760 = n5825 & n1759 ;
  assign n5826 = ~n1754 ;
  assign n1761 = n1749 & n5826 ;
  assign n1762 = n1755 | n1761 ;
  assign n5827 = ~n1762 ;
  assign n1764 = n1760 & n5827 ;
  assign n1765 = n1755 | n1764 ;
  assign n1767 = n1744 & n1765 ;
  assign n5828 = ~n1765 ;
  assign n1766 = n1744 & n5828 ;
  assign n5829 = ~n1744 ;
  assign n1768 = n5829 & n1765 ;
  assign n1769 = n1766 | n1768 ;
  assign n1645 = n1642 | n1644 ;
  assign n5830 = ~n1646 ;
  assign n1770 = n1645 & n5830 ;
  assign n1772 = n1769 & n1770 ;
  assign n1773 = n1767 | n1772 ;
  assign n5831 = ~n1647 ;
  assign n1650 = n5831 & n1649 ;
  assign n5832 = ~n1649 ;
  assign n1774 = n1647 & n5832 ;
  assign n1775 = n1650 | n1774 ;
  assign n1776 = n1773 & n1775 ;
  assign n1701 = n1698 | n1700 ;
  assign n1777 = n1698 & n1700 ;
  assign n5833 = ~n1777 ;
  assign n1778 = n1701 & n5833 ;
  assign n1779 = n1773 | n1775 ;
  assign n5834 = ~n1776 ;
  assign n1780 = n5834 & n1779 ;
  assign n5835 = ~n1778 ;
  assign n1782 = n5835 & n1780 ;
  assign n1783 = n1776 | n1782 ;
  assign n5836 = ~n1709 ;
  assign n1784 = n5836 & n1710 ;
  assign n1785 = n1711 | n1784 ;
  assign n5837 = ~n1785 ;
  assign n1786 = n1783 & n5837 ;
  assign n1787 = n545 | n1618 ;
  assign n1431 = n859 & n1428 ;
  assign n1375 = n5554 & n1373 ;
  assign n1788 = n851 & n1385 ;
  assign n1789 = n1375 | n1788 ;
  assign n1790 = n5512 & n1434 ;
  assign n5838 = ~n1790 ;
  assign n1791 = n1789 & n5838 ;
  assign n5839 = ~n1431 ;
  assign n1792 = n5839 & n1791 ;
  assign n1233 = n1064 & n1229 ;
  assign n1083 = n5721 & n891 ;
  assign n1793 = n274 & n893 ;
  assign n1794 = n1083 | n1793 ;
  assign n1795 = n895 & n5722 ;
  assign n5840 = ~n1795 ;
  assign n1796 = n1794 & n5840 ;
  assign n5841 = ~n1233 ;
  assign n1797 = n5841 & n1796 ;
  assign n1798 = n1792 & n1797 ;
  assign n1271 = n1052 | n1265 ;
  assign n1260 = n5647 & n1251 ;
  assign n1799 = n1043 & n1264 ;
  assign n1800 = n1260 | n1799 ;
  assign n5842 = ~n1800 ;
  assign n1801 = n1271 & n5842 ;
  assign n1802 = n1052 & n1324 ;
  assign n5843 = ~n1802 ;
  assign n1803 = n1801 & n5843 ;
  assign n1804 = n1792 | n1797 ;
  assign n5844 = ~n1798 ;
  assign n1805 = n5844 & n1804 ;
  assign n1807 = n1803 & n1805 ;
  assign n1808 = n1798 | n1807 ;
  assign n1809 = n5797 & n1808 ;
  assign n1810 = n1787 & n1809 ;
  assign n5845 = ~n1810 ;
  assign n1812 = n1808 & n5845 ;
  assign n1811 = n1619 | n1810 ;
  assign n5846 = ~n1811 ;
  assign n1813 = n1787 & n5846 ;
  assign n1814 = n1812 | n1813 ;
  assign n1741 = n1727 | n1740 ;
  assign n5847 = ~n1743 ;
  assign n1815 = n1741 & n5847 ;
  assign n1816 = n1814 & n1815 ;
  assign n1817 = n1810 | n1816 ;
  assign n5848 = ~n1691 ;
  assign n1692 = n1686 & n5848 ;
  assign n5849 = ~n1687 ;
  assign n1818 = n1686 & n5849 ;
  assign n1819 = n1689 | n1818 ;
  assign n5850 = ~n1692 ;
  assign n1820 = n5850 & n1819 ;
  assign n5851 = ~n1820 ;
  assign n1822 = n1817 & n5851 ;
  assign n5852 = ~n1817 ;
  assign n1821 = n5852 & n1820 ;
  assign n1823 = n1821 | n1822 ;
  assign n1771 = n1769 | n1770 ;
  assign n5853 = ~n1772 ;
  assign n1824 = n1771 & n5853 ;
  assign n5854 = ~n1823 ;
  assign n1826 = n5854 & n1824 ;
  assign n1827 = n1822 | n1826 ;
  assign n1781 = n1778 & n1780 ;
  assign n1828 = n1778 | n1780 ;
  assign n5855 = ~n1781 ;
  assign n1829 = n5855 & n1828 ;
  assign n5856 = ~n1829 ;
  assign n1830 = n1827 & n5856 ;
  assign n1607 = n672 & n5765 ;
  assign n1832 = n5514 & n1545 ;
  assign n1831 = n859 | n1177 ;
  assign n1833 = n1544 & n1831 ;
  assign n1834 = n1832 | n1833 ;
  assign n1835 = n1607 | n1834 ;
  assign n1436 = n5554 & n1434 ;
  assign n1380 = n1052 | n1373 ;
  assign n1836 = n1052 & n5675 ;
  assign n5857 = ~n1836 ;
  assign n1837 = n1380 & n5857 ;
  assign n5858 = ~n1436 ;
  assign n1838 = n5858 & n1837 ;
  assign n1839 = n851 & n1428 ;
  assign n5859 = ~n1839 ;
  assign n1840 = n1838 & n5859 ;
  assign n5860 = ~n1835 ;
  assign n1842 = n5860 & n1840 ;
  assign n1267 = n1043 | n1265 ;
  assign n1261 = n5722 & n1251 ;
  assign n1843 = n1229 & n1264 ;
  assign n1844 = n1261 | n1843 ;
  assign n5861 = ~n1844 ;
  assign n1845 = n1267 & n5861 ;
  assign n1846 = n1043 & n1324 ;
  assign n5862 = ~n1846 ;
  assign n1847 = n1845 & n5862 ;
  assign n1841 = n1835 | n1840 ;
  assign n1848 = n1835 & n1840 ;
  assign n5863 = ~n1848 ;
  assign n1849 = n1841 & n5863 ;
  assign n5864 = ~n1849 ;
  assign n1851 = n1847 & n5864 ;
  assign n1852 = n1842 | n1851 ;
  assign n877 = n275 & n868 ;
  assign n714 = n5499 & n708 ;
  assign n1853 = n282 & n716 ;
  assign n1854 = n714 | n1853 ;
  assign n1855 = n5498 & n717 ;
  assign n5865 = ~n1855 ;
  assign n1856 = n1854 & n5865 ;
  assign n5866 = ~n877 ;
  assign n1857 = n5866 & n1856 ;
  assign n1726 = n1721 | n1725 ;
  assign n1858 = n1721 & n1725 ;
  assign n5867 = ~n1858 ;
  assign n1859 = n1726 & n5867 ;
  assign n1860 = n1857 & n1859 ;
  assign n1861 = n1857 | n1859 ;
  assign n5868 = ~n1860 ;
  assign n1862 = n5868 & n1861 ;
  assign n5869 = ~n1862 ;
  assign n1864 = n1852 & n5869 ;
  assign n5870 = ~n1859 ;
  assign n1865 = n1857 & n5870 ;
  assign n1866 = n1864 | n1865 ;
  assign n1763 = n1760 & n1762 ;
  assign n1867 = n1760 | n1762 ;
  assign n5871 = ~n1763 ;
  assign n1868 = n5871 & n1867 ;
  assign n5872 = ~n1868 ;
  assign n1870 = n1866 & n5872 ;
  assign n1871 = n1814 | n1815 ;
  assign n5873 = ~n1816 ;
  assign n1872 = n5873 & n1871 ;
  assign n5874 = ~n1866 ;
  assign n1869 = n5874 & n1868 ;
  assign n1873 = n1869 | n1870 ;
  assign n5875 = ~n1873 ;
  assign n1875 = n1872 & n5875 ;
  assign n1876 = n1870 | n1875 ;
  assign n1437 = n5595 & n1434 ;
  assign n1381 = n1043 | n1373 ;
  assign n1908 = n1043 & n5675 ;
  assign n5876 = ~n1908 ;
  assign n1909 = n1381 & n5876 ;
  assign n5877 = ~n1437 ;
  assign n1910 = n5877 & n1909 ;
  assign n1911 = n1052 & n1428 ;
  assign n5878 = ~n1911 ;
  assign n1912 = n1910 & n5878 ;
  assign n1269 = n1229 | n1265 ;
  assign n1262 = n5721 & n1251 ;
  assign n1913 = n274 & n1264 ;
  assign n1914 = n1262 | n1913 ;
  assign n5879 = ~n1914 ;
  assign n1915 = n1269 & n5879 ;
  assign n1916 = n1229 & n1324 ;
  assign n5880 = ~n1916 ;
  assign n1917 = n1915 & n5880 ;
  assign n1924 = n1912 & n1917 ;
  assign n1070 = n275 & n1064 ;
  assign n1084 = n5499 & n891 ;
  assign n1919 = n282 & n893 ;
  assign n1920 = n1084 | n1919 ;
  assign n1921 = n5498 & n895 ;
  assign n5881 = ~n1921 ;
  assign n1922 = n1920 & n5881 ;
  assign n5882 = ~n1070 ;
  assign n1923 = n5882 & n1922 ;
  assign n1918 = n1912 | n1917 ;
  assign n5883 = ~n1924 ;
  assign n1925 = n1918 & n5883 ;
  assign n1927 = n1923 & n1925 ;
  assign n1928 = n1924 | n1927 ;
  assign n5884 = ~n1847 ;
  assign n1850 = n5884 & n1849 ;
  assign n1929 = n1850 | n1851 ;
  assign n5885 = ~n1929 ;
  assign n1931 = n1928 & n5885 ;
  assign n1074 = n274 & n1064 ;
  assign n1076 = n5498 & n891 ;
  assign n1877 = n275 & n893 ;
  assign n1878 = n1076 | n1877 ;
  assign n1879 = n5721 & n895 ;
  assign n5886 = ~n1879 ;
  assign n1880 = n1878 & n5886 ;
  assign n5887 = ~n1074 ;
  assign n1881 = n5887 & n1880 ;
  assign n1608 = n859 & n5765 ;
  assign n1883 = n5512 & n1545 ;
  assign n1882 = n851 | n1177 ;
  assign n1884 = n1544 & n1882 ;
  assign n1885 = n1883 | n1884 ;
  assign n1886 = n1608 | n1885 ;
  assign n1887 = n282 & n890 ;
  assign n1888 = n846 | n1887 ;
  assign n1889 = n282 & n1064 ;
  assign n5888 = ~n1889 ;
  assign n1890 = n1888 & n5888 ;
  assign n1892 = n846 & n1890 ;
  assign n5889 = ~n1886 ;
  assign n1894 = n5889 & n1892 ;
  assign n1895 = n1881 & n1894 ;
  assign n1896 = n1881 | n1894 ;
  assign n5890 = ~n1895 ;
  assign n1897 = n5890 & n1896 ;
  assign n5891 = ~n1897 ;
  assign n1898 = n1722 & n5891 ;
  assign n5892 = ~n1722 ;
  assign n1932 = n5892 & n1897 ;
  assign n1933 = n1898 | n1932 ;
  assign n1930 = n1928 & n1929 ;
  assign n1934 = n1928 | n1929 ;
  assign n5893 = ~n1930 ;
  assign n1935 = n5893 & n1934 ;
  assign n5894 = ~n1935 ;
  assign n1937 = n1933 & n5894 ;
  assign n1938 = n1931 | n1937 ;
  assign n1891 = n846 | n1890 ;
  assign n1939 = n1052 & n5765 ;
  assign n1941 = n5595 & n1545 ;
  assign n1940 = n1043 | n1177 ;
  assign n1942 = n1544 & n1940 ;
  assign n1943 = n1941 | n1942 ;
  assign n1944 = n1939 | n1943 ;
  assign n1945 = n282 & n5651 ;
  assign n1946 = n1037 | n1945 ;
  assign n1947 = n282 & n1324 ;
  assign n5895 = ~n1947 ;
  assign n1948 = n1946 & n5895 ;
  assign n1949 = n1037 & n1948 ;
  assign n5896 = ~n1944 ;
  assign n1951 = n5896 & n1949 ;
  assign n5897 = ~n1892 ;
  assign n1952 = n5897 & n1951 ;
  assign n1954 = n1891 & n1952 ;
  assign n1438 = n5722 & n1434 ;
  assign n1382 = n274 | n1373 ;
  assign n1956 = n274 & n5675 ;
  assign n5898 = ~n1956 ;
  assign n1957 = n1382 & n5898 ;
  assign n5899 = ~n1438 ;
  assign n1958 = n5899 & n1957 ;
  assign n1959 = n1229 & n1428 ;
  assign n5900 = ~n1959 ;
  assign n1960 = n1958 & n5900 ;
  assign n1273 = n275 | n1265 ;
  assign n1256 = n5499 & n1251 ;
  assign n1961 = n282 & n1264 ;
  assign n1962 = n1256 | n1961 ;
  assign n5901 = ~n1962 ;
  assign n1963 = n1273 & n5901 ;
  assign n1964 = n275 & n1324 ;
  assign n5902 = ~n1964 ;
  assign n1965 = n1963 & n5902 ;
  assign n1967 = n1960 & n1965 ;
  assign n1966 = n1960 | n1965 ;
  assign n1950 = n1944 & n1949 ;
  assign n1968 = n1944 | n1949 ;
  assign n5903 = ~n1950 ;
  assign n1969 = n5903 & n1968 ;
  assign n5904 = ~n1969 ;
  assign n1970 = n1966 & n5904 ;
  assign n1971 = n1967 | n1970 ;
  assign n5905 = ~n1954 ;
  assign n1955 = n1951 & n5905 ;
  assign n1953 = n1891 & n1951 ;
  assign n1972 = n1892 | n1953 ;
  assign n5906 = ~n1972 ;
  assign n1973 = n1891 & n5906 ;
  assign n1974 = n1955 | n1973 ;
  assign n1976 = n1971 & n1974 ;
  assign n1977 = n1954 | n1976 ;
  assign n1327 = n274 & n1324 ;
  assign n1254 = n275 | n1251 ;
  assign n1978 = n275 & n5702 ;
  assign n5907 = ~n1978 ;
  assign n1979 = n1254 & n5907 ;
  assign n1980 = n274 | n1265 ;
  assign n5908 = ~n1979 ;
  assign n1981 = n5908 & n1980 ;
  assign n5909 = ~n1327 ;
  assign n1982 = n5909 & n1981 ;
  assign n1432 = n1043 & n1428 ;
  assign n1378 = n5722 & n1373 ;
  assign n1983 = n1229 & n1385 ;
  assign n1984 = n1378 | n1983 ;
  assign n1985 = n5647 & n1434 ;
  assign n5910 = ~n1985 ;
  assign n1986 = n1984 & n5910 ;
  assign n5911 = ~n1432 ;
  assign n1987 = n5911 & n1986 ;
  assign n1609 = n851 & n5765 ;
  assign n1989 = n5554 & n1545 ;
  assign n1988 = n1052 | n1177 ;
  assign n1990 = n1544 & n1988 ;
  assign n1991 = n1989 | n1990 ;
  assign n1992 = n1609 | n1991 ;
  assign n5912 = ~n1992 ;
  assign n1993 = n1987 & n5912 ;
  assign n5913 = ~n1987 ;
  assign n1994 = n5913 & n1992 ;
  assign n1995 = n1993 | n1994 ;
  assign n5914 = ~n1982 ;
  assign n1996 = n5914 & n1995 ;
  assign n5915 = ~n1995 ;
  assign n1997 = n1982 & n5915 ;
  assign n1611 = n1043 & n5765 ;
  assign n1999 = n5647 & n1545 ;
  assign n1998 = n1177 | n1229 ;
  assign n2000 = n1544 & n1998 ;
  assign n2001 = n1999 | n2000 ;
  assign n2002 = n1611 | n2001 ;
  assign n1439 = n5721 & n1434 ;
  assign n1383 = n275 | n1373 ;
  assign n2003 = n275 & n5675 ;
  assign n5916 = ~n2003 ;
  assign n2004 = n1383 & n5916 ;
  assign n5917 = ~n1439 ;
  assign n2005 = n5917 & n2004 ;
  assign n2006 = n274 & n1428 ;
  assign n5918 = ~n2006 ;
  assign n2007 = n2005 & n5918 ;
  assign n2008 = n2002 | n2007 ;
  assign n2009 = n2002 & n2007 ;
  assign n5919 = ~n2009 ;
  assign n2010 = n2008 & n5919 ;
  assign n1610 = n1229 & n5765 ;
  assign n2012 = n5722 & n1545 ;
  assign n2011 = n274 | n1177 ;
  assign n2013 = n1544 & n2011 ;
  assign n2014 = n2012 | n2013 ;
  assign n2015 = n1610 | n2014 ;
  assign n2016 = n282 & n1372 ;
  assign n2017 = n1227 | n2016 ;
  assign n2018 = n282 & n1428 ;
  assign n5920 = ~n2018 ;
  assign n2019 = n2017 & n5920 ;
  assign n2021 = n1227 & n2019 ;
  assign n5921 = ~n2015 ;
  assign n2022 = n5921 & n2021 ;
  assign n5922 = ~n2022 ;
  assign n2023 = n2010 & n5922 ;
  assign n5923 = ~n2010 ;
  assign n2024 = n5923 & n2022 ;
  assign n2026 = n274 & n5765 ;
  assign n2027 = n5721 & n1545 ;
  assign n1178 = n275 | n1177 ;
  assign n2028 = n1178 & n1544 ;
  assign n2029 = n2027 | n2028 ;
  assign n2030 = n2026 | n2029 ;
  assign n1546 = n275 & n5766 ;
  assign n2031 = n282 | n1177 ;
  assign n2032 = n1546 | n2031 ;
  assign n2033 = n2030 | n2032 ;
  assign n2020 = n1227 | n2019 ;
  assign n2034 = n2030 & n2032 ;
  assign n2035 = n2021 | n2034 ;
  assign n5924 = ~n2035 ;
  assign n2036 = n2020 & n5924 ;
  assign n5925 = ~n2036 ;
  assign n2037 = n2033 & n5925 ;
  assign n5926 = ~n2021 ;
  assign n2038 = n2015 & n5926 ;
  assign n2039 = n2022 | n2038 ;
  assign n2040 = n2037 | n2039 ;
  assign n2025 = n275 & n1428 ;
  assign n1440 = n5498 & n1434 ;
  assign n2041 = n282 & n5675 ;
  assign n2042 = n282 | n1373 ;
  assign n2043 = n2037 & n2039 ;
  assign n5927 = ~n2043 ;
  assign n2044 = n2042 & n5927 ;
  assign n5928 = ~n2041 ;
  assign n2045 = n5928 & n2044 ;
  assign n5929 = ~n1440 ;
  assign n2046 = n5929 & n2045 ;
  assign n5930 = ~n2025 ;
  assign n2047 = n5930 & n2046 ;
  assign n5931 = ~n2047 ;
  assign n2048 = n2040 & n5931 ;
  assign n5932 = ~n1945 ;
  assign n2049 = n5932 & n2048 ;
  assign n2050 = n2024 | n2049 ;
  assign n2051 = n2023 | n2050 ;
  assign n5933 = ~n2048 ;
  assign n2052 = n1945 & n5933 ;
  assign n5934 = ~n2052 ;
  assign n2053 = n2051 & n5934 ;
  assign n5935 = ~n1949 ;
  assign n2054 = n1944 & n5935 ;
  assign n2055 = n1951 | n2054 ;
  assign n5936 = ~n1967 ;
  assign n2057 = n1966 & n5936 ;
  assign n2058 = n2055 | n2057 ;
  assign n5937 = ~n2055 ;
  assign n2056 = n1966 & n5937 ;
  assign n2059 = n1967 | n2056 ;
  assign n5938 = ~n2059 ;
  assign n2060 = n1966 & n5938 ;
  assign n5939 = ~n2060 ;
  assign n2061 = n2058 & n5939 ;
  assign n2062 = n2053 & n2061 ;
  assign n5940 = ~n2002 ;
  assign n2063 = n5940 & n2007 ;
  assign n2064 = n2024 | n2063 ;
  assign n5941 = ~n2062 ;
  assign n2065 = n5941 & n2064 ;
  assign n2066 = n2053 | n2061 ;
  assign n5942 = ~n2065 ;
  assign n2067 = n5942 & n2066 ;
  assign n5943 = ~n1974 ;
  assign n1975 = n1971 & n5943 ;
  assign n5944 = ~n1971 ;
  assign n2068 = n5944 & n1974 ;
  assign n2069 = n1975 | n2068 ;
  assign n5945 = ~n2069 ;
  assign n2070 = n2067 & n5945 ;
  assign n2071 = n1997 | n2070 ;
  assign n2072 = n1996 | n2071 ;
  assign n5946 = ~n2067 ;
  assign n2073 = n5946 & n2069 ;
  assign n5947 = ~n2073 ;
  assign n2074 = n2072 & n5947 ;
  assign n5948 = ~n2074 ;
  assign n2076 = n1977 & n5948 ;
  assign n5949 = ~n1977 ;
  assign n2075 = n5949 & n2074 ;
  assign n5950 = ~n1925 ;
  assign n1926 = n1923 & n5950 ;
  assign n5951 = ~n1923 ;
  assign n2077 = n5951 & n1925 ;
  assign n2078 = n1926 | n2077 ;
  assign n1893 = n1886 | n1892 ;
  assign n2079 = n1886 & n1892 ;
  assign n5952 = ~n2079 ;
  assign n2080 = n1893 & n5952 ;
  assign n2081 = n1993 | n1997 ;
  assign n5953 = ~n2081 ;
  assign n2082 = n2080 & n5953 ;
  assign n5954 = ~n2080 ;
  assign n2083 = n5954 & n2081 ;
  assign n2084 = n2082 | n2083 ;
  assign n2085 = n2078 | n2084 ;
  assign n2086 = n2078 & n2084 ;
  assign n5955 = ~n2086 ;
  assign n2087 = n2085 & n5955 ;
  assign n2088 = n2075 | n2087 ;
  assign n5956 = ~n2076 ;
  assign n2089 = n5956 & n2088 ;
  assign n5957 = ~n2084 ;
  assign n2090 = n2078 & n5957 ;
  assign n2091 = n2083 | n2090 ;
  assign n5958 = ~n2089 ;
  assign n2093 = n5958 & n2091 ;
  assign n5959 = ~n2091 ;
  assign n2092 = n2089 & n5959 ;
  assign n1936 = n1933 & n1935 ;
  assign n2094 = n1933 | n1935 ;
  assign n5960 = ~n1936 ;
  assign n2095 = n5960 & n2094 ;
  assign n2096 = n2092 | n2095 ;
  assign n5961 = ~n2093 ;
  assign n2097 = n5961 & n2096 ;
  assign n5962 = ~n2097 ;
  assign n2098 = n1938 & n5962 ;
  assign n1899 = n1722 & n1897 ;
  assign n1900 = n1895 | n1899 ;
  assign n1806 = n1803 | n1805 ;
  assign n5963 = ~n1807 ;
  assign n1901 = n1806 & n5963 ;
  assign n5964 = ~n1900 ;
  assign n1902 = n5964 & n1901 ;
  assign n5965 = ~n1901 ;
  assign n1903 = n1900 & n5965 ;
  assign n1904 = n1902 | n1903 ;
  assign n1863 = n1852 & n1862 ;
  assign n1905 = n1852 | n1862 ;
  assign n5966 = ~n1863 ;
  assign n1906 = n5966 & n1905 ;
  assign n5967 = ~n1904 ;
  assign n1907 = n5967 & n1906 ;
  assign n5968 = ~n1906 ;
  assign n2099 = n1904 & n5968 ;
  assign n5969 = ~n1938 ;
  assign n2100 = n5969 & n2097 ;
  assign n2101 = n2099 | n2100 ;
  assign n2102 = n1907 | n2101 ;
  assign n5970 = ~n2098 ;
  assign n2103 = n5970 & n2102 ;
  assign n2104 = n1900 & n1901 ;
  assign n2105 = n2099 | n2104 ;
  assign n5971 = ~n2103 ;
  assign n2107 = n5971 & n2105 ;
  assign n5972 = ~n2105 ;
  assign n2106 = n2103 & n5972 ;
  assign n1874 = n1872 & n1873 ;
  assign n2108 = n1872 | n1873 ;
  assign n5973 = ~n1874 ;
  assign n2109 = n5973 & n2108 ;
  assign n2110 = n2106 | n2109 ;
  assign n5974 = ~n2107 ;
  assign n2111 = n5974 & n2110 ;
  assign n5975 = ~n2111 ;
  assign n2112 = n1876 & n5975 ;
  assign n5976 = ~n1824 ;
  assign n1825 = n1823 & n5976 ;
  assign n5977 = ~n1876 ;
  assign n2113 = n5977 & n2111 ;
  assign n2114 = n1825 | n2113 ;
  assign n2115 = n1826 | n2114 ;
  assign n5978 = ~n2112 ;
  assign n2116 = n5978 & n2115 ;
  assign n5979 = ~n1827 ;
  assign n2117 = n5979 & n1829 ;
  assign n2118 = n2116 | n2117 ;
  assign n5980 = ~n1830 ;
  assign n2119 = n5980 & n2118 ;
  assign n5981 = ~n1783 ;
  assign n2120 = n5981 & n1785 ;
  assign n2121 = n1786 | n2120 ;
  assign n2122 = n2119 | n2121 ;
  assign n5982 = ~n1786 ;
  assign n2123 = n5982 & n2122 ;
  assign n1715 = n1712 | n1714 ;
  assign n2124 = n1712 & n1714 ;
  assign n5983 = ~n2124 ;
  assign n2125 = n1715 & n5983 ;
  assign n2127 = n2123 | n2125 ;
  assign n5984 = ~n1716 ;
  assign n2128 = n5984 & n2127 ;
  assign n1674 = n1671 | n1673 ;
  assign n2129 = n1671 & n1673 ;
  assign n5985 = ~n2129 ;
  assign n2130 = n1674 & n5985 ;
  assign n2131 = n2128 | n2130 ;
  assign n5986 = ~n1675 ;
  assign n2132 = n5986 & n2131 ;
  assign n2134 = n1602 | n2132 ;
  assign n5987 = ~n1601 ;
  assign n2135 = n5987 & n2134 ;
  assign n5988 = ~n1487 ;
  assign n1490 = n5988 & n1489 ;
  assign n2136 = n1490 | n1491 ;
  assign n2137 = n2135 | n2136 ;
  assign n5989 = ~n1491 ;
  assign n2138 = n5989 & n2137 ;
  assign n2140 = n1360 | n2138 ;
  assign n5990 = ~n1359 ;
  assign n2141 = n5990 & n2140 ;
  assign n1309 = n1306 | n1308 ;
  assign n2142 = n1306 & n1308 ;
  assign n5991 = ~n2142 ;
  assign n2143 = n1309 & n5991 ;
  assign n2144 = n2141 | n2143 ;
  assign n5992 = ~n1310 ;
  assign n2145 = n5992 & n2144 ;
  assign n2147 = n1125 | n2145 ;
  assign n5993 = ~n1124 ;
  assign n2148 = n5993 & n2147 ;
  assign n915 = n867 & n913 ;
  assign n5994 = ~n919 ;
  assign n921 = n917 & n5994 ;
  assign n922 = n915 | n921 ;
  assign n686 = n523 & n685 ;
  assign n695 = n5540 & n694 ;
  assign n701 = n528 & n543 ;
  assign n702 = n695 | n701 ;
  assign n703 = n5542 & n692 ;
  assign n5995 = ~n703 ;
  assign n704 = n702 & n5995 ;
  assign n5996 = ~n686 ;
  assign n705 = n5996 & n704 ;
  assign n730 = n722 | n729 ;
  assign n5997 = ~n730 ;
  assign n731 = n705 & n5997 ;
  assign n5998 = ~n705 ;
  assign n733 = n5998 & n730 ;
  assign n734 = n731 | n733 ;
  assign n674 = n5549 & n673 ;
  assign n675 = n666 & n5587 ;
  assign n676 = n674 | n675 ;
  assign n678 = n441 & n677 ;
  assign n5999 = ~n676 ;
  assign n679 = n5999 & n678 ;
  assign n6000 = ~n678 ;
  assign n735 = n676 & n6000 ;
  assign n736 = n679 | n735 ;
  assign n6001 = ~n736 ;
  assign n737 = n734 & n6001 ;
  assign n6002 = ~n734 ;
  assign n923 = n6002 & n736 ;
  assign n924 = n737 | n923 ;
  assign n925 = n922 | n924 ;
  assign n2149 = n922 & n924 ;
  assign n6003 = ~n2149 ;
  assign n2150 = n925 & n6003 ;
  assign n2151 = n2148 | n2150 ;
  assign n2227 = n2148 & n2150 ;
  assign n6004 = ~n2227 ;
  assign n2228 = n2151 & n6004 ;
  assign n6005 = ~n2228 ;
  assign n2229 = n2226 & n6005 ;
  assign n6006 = ~n2226 ;
  assign n2230 = n6006 & n2228 ;
  assign n2166 = n131 | n467 ;
  assign n2167 = n217 | n2166 ;
  assign n327 = n325 | n326 ;
  assign n328 = n253 | n327 ;
  assign n2183 = n358 | n994 ;
  assign n2184 = n139 | n2183 ;
  assign n2232 = n328 | n2184 ;
  assign n2233 = n234 | n2232 ;
  assign n2234 = n298 | n2233 ;
  assign n2235 = n636 | n2234 ;
  assign n2236 = n2167 | n2235 ;
  assign n2237 = n352 | n2236 ;
  assign n2238 = n219 | n2237 ;
  assign n2239 = n391 | n2238 ;
  assign n2240 = n223 | n2239 ;
  assign n2241 = n204 | n2240 ;
  assign n2242 = n252 | n932 ;
  assign n2243 = n446 | n2242 ;
  assign n2244 = n145 | n2243 ;
  assign n2245 = n108 | n2244 ;
  assign n2246 = n236 | n2245 ;
  assign n2247 = n580 | n627 ;
  assign n2248 = n2246 | n2247 ;
  assign n2249 = n225 | n2248 ;
  assign n2250 = n414 | n2249 ;
  assign n2251 = n120 | n2250 ;
  assign n2252 = n752 | n2251 ;
  assign n2253 = n175 | n505 ;
  assign n2254 = n470 | n2253 ;
  assign n2255 = n299 | n310 ;
  assign n2256 = n444 | n2255 ;
  assign n2257 = n477 | n2256 ;
  assign n2258 = n2254 | n2257 ;
  assign n2259 = n153 | n2258 ;
  assign n2260 = n576 | n2259 ;
  assign n2261 = n643 | n2260 ;
  assign n2262 = n2252 | n2261 ;
  assign n2263 = n2241 | n2262 ;
  assign n2264 = n314 | n2263 ;
  assign n2265 = n333 | n2264 ;
  assign n2266 = n553 | n2265 ;
  assign n2146 = n1125 & n2145 ;
  assign n6007 = ~n2146 ;
  assign n2267 = n6007 & n2147 ;
  assign n6008 = ~n2267 ;
  assign n2269 = n2266 & n6008 ;
  assign n2270 = n393 | n2254 ;
  assign n2271 = n450 | n2270 ;
  assign n2272 = n136 | n2271 ;
  assign n2273 = n186 | n2272 ;
  assign n2274 = n126 | n2273 ;
  assign n2275 = n356 | n2274 ;
  assign n2276 = n332 | n2275 ;
  assign n2277 = n364 | n2276 ;
  assign n2278 = n598 | n2277 ;
  assign n2192 = n137 | n808 ;
  assign n2193 = n296 | n2192 ;
  assign n2194 = n457 | n2193 ;
  assign n2195 = n354 | n2194 ;
  assign n2196 = n145 | n2195 ;
  assign n2197 = n552 | n2196 ;
  assign n2279 = n446 | n551 ;
  assign n2280 = n235 | n2279 ;
  assign n2281 = n149 | n2241 ;
  assign n2282 = n293 | n2281 ;
  assign n2283 = n213 | n2282 ;
  assign n2284 = n1516 | n2283 ;
  assign n2285 = n2280 | n2284 ;
  assign n6009 = ~n2285 ;
  assign n2286 = n322 & n6009 ;
  assign n6010 = ~n2197 ;
  assign n2287 = n6010 & n2286 ;
  assign n6011 = ~n2278 ;
  assign n2288 = n6011 & n2287 ;
  assign n6012 = ~n1006 ;
  assign n2289 = n6012 & n2288 ;
  assign n6013 = ~n173 ;
  assign n2290 = n6013 & n2289 ;
  assign n6014 = ~n340 ;
  assign n2291 = n6014 & n2290 ;
  assign n2292 = n5611 & n2291 ;
  assign n2293 = n5725 & n2292 ;
  assign n6015 = ~n310 ;
  assign n2294 = n6015 & n2293 ;
  assign n2295 = n2141 & n2143 ;
  assign n6016 = ~n2295 ;
  assign n2296 = n2144 & n6016 ;
  assign n2298 = n2294 | n2296 ;
  assign n2297 = n2294 & n2296 ;
  assign n2300 = n135 | n225 ;
  assign n2301 = n120 | n2300 ;
  assign n2302 = n169 | n2301 ;
  assign n2303 = n232 | n2302 ;
  assign n2304 = n354 | n2303 ;
  assign n2305 = n214 | n2304 ;
  assign n2306 = n165 | n2305 ;
  assign n366 = n124 | n365 ;
  assign n2307 = n138 | n1163 ;
  assign n2308 = n970 | n2307 ;
  assign n2309 = n643 | n2308 ;
  assign n2310 = n366 | n2309 ;
  assign n2311 = n334 | n2310 ;
  assign n2312 = n457 | n2311 ;
  assign n2313 = n446 | n2312 ;
  assign n2314 = n344 | n2313 ;
  assign n2315 = n101 | n949 ;
  assign n2316 = n323 | n2315 ;
  assign n2317 = n215 | n226 ;
  assign n2318 = n143 | n2317 ;
  assign n2319 = n209 | n2318 ;
  assign n2320 = n468 | n2319 ;
  assign n2321 = n2316 | n2320 ;
  assign n2322 = n2314 | n2321 ;
  assign n2323 = n2306 | n2322 ;
  assign n2324 = n325 | n2323 ;
  assign n2325 = n405 | n2324 ;
  assign n2326 = n192 | n2325 ;
  assign n2327 = n217 | n2326 ;
  assign n2328 = n295 | n2327 ;
  assign n2329 = n449 | n2328 ;
  assign n2330 = n444 | n2329 ;
  assign n2139 = n1360 & n2138 ;
  assign n6017 = ~n2139 ;
  assign n2331 = n6017 & n2140 ;
  assign n6018 = ~n2331 ;
  assign n2333 = n2330 & n6018 ;
  assign n2334 = n211 | n507 ;
  assign n2335 = n752 | n2334 ;
  assign n2336 = n342 | n2335 ;
  assign n2337 = n300 | n775 ;
  assign n2338 = n957 | n2337 ;
  assign n2339 = n166 | n2338 ;
  assign n2340 = n110 | n2339 ;
  assign n2341 = n323 | n2340 ;
  assign n2342 = n468 | n2341 ;
  assign n2343 = n135 | n143 ;
  assign n2344 = n101 | n345 ;
  assign n2345 = n236 | n2344 ;
  assign n2346 = n429 | n2345 ;
  assign n2347 = n2343 | n2346 ;
  assign n2348 = n1153 | n2347 ;
  assign n2349 = n341 | n2348 ;
  assign n2350 = n311 | n2349 ;
  assign n2351 = n2342 | n2350 ;
  assign n2352 = n1021 | n2351 ;
  assign n2353 = n956 | n2352 ;
  assign n2354 = n2336 | n2353 ;
  assign n2355 = n149 | n2354 ;
  assign n2356 = n215 | n2355 ;
  assign n2357 = n494 | n2356 ;
  assign n2358 = n2135 & n2136 ;
  assign n6019 = ~n2358 ;
  assign n2359 = n2137 & n6019 ;
  assign n6020 = ~n2359 ;
  assign n2360 = n2357 & n6020 ;
  assign n6021 = ~n2357 ;
  assign n2361 = n6021 & n2359 ;
  assign n2363 = n138 | n309 ;
  assign n2364 = n414 | n2363 ;
  assign n2365 = n310 | n2364 ;
  assign n2366 = n222 | n2365 ;
  assign n2367 = n552 | n2366 ;
  assign n2368 = n233 | n2367 ;
  assign n2369 = n253 | n448 ;
  assign n2370 = n553 | n2369 ;
  assign n2371 = n192 | n235 ;
  assign n2372 = n2370 | n2371 ;
  assign n2373 = n936 | n2372 ;
  assign n2374 = n186 | n2373 ;
  assign n2375 = n324 | n2374 ;
  assign n2376 = n345 | n2375 ;
  assign n2377 = n326 | n2376 ;
  assign n2378 = n189 | n2377 ;
  assign n2379 = n502 | n2378 ;
  assign n368 = n366 | n367 ;
  assign n369 = n364 | n368 ;
  assign n371 = n369 | n370 ;
  assign n372 = n363 | n371 ;
  assign n373 = n352 | n372 ;
  assign n374 = n171 | n373 ;
  assign n375 = n130 | n374 ;
  assign n376 = n143 | n375 ;
  assign n377 = n221 | n376 ;
  assign n378 = n153 | n377 ;
  assign n379 = n347 | n378 ;
  assign n2380 = n379 | n447 ;
  assign n2381 = n2379 | n2380 ;
  assign n2382 = n769 | n2381 ;
  assign n2383 = n2368 | n2382 ;
  assign n2384 = n194 | n2383 ;
  assign n2385 = n219 | n2384 ;
  assign n2386 = n391 | n2385 ;
  assign n2387 = n164 | n2386 ;
  assign n2388 = n344 | n2387 ;
  assign n2389 = n471 | n2388 ;
  assign n2133 = n1602 & n2132 ;
  assign n6022 = ~n2133 ;
  assign n2390 = n6022 & n2134 ;
  assign n6023 = ~n2390 ;
  assign n2392 = n2389 & n6023 ;
  assign n2393 = n563 | n2256 ;
  assign n2394 = n932 | n2393 ;
  assign n2395 = n408 | n2394 ;
  assign n2396 = n357 | n2395 ;
  assign n2397 = n110 | n2396 ;
  assign n2398 = n323 | n2397 ;
  assign n2399 = n221 | n2398 ;
  assign n2400 = n413 | n472 ;
  assign n2401 = n295 | n2400 ;
  assign n2402 = n114 | n2401 ;
  assign n2403 = n222 | n2402 ;
  assign n2404 = n364 | n2403 ;
  assign n2405 = n589 | n2404 ;
  assign n2406 = n2399 | n2405 ;
  assign n2407 = n768 | n2406 ;
  assign n2408 = n1012 | n2407 ;
  assign n2409 = n146 | n2408 ;
  assign n2410 = n226 | n2409 ;
  assign n2411 = n217 | n2410 ;
  assign n2412 = n224 | n2411 ;
  assign n2413 = n333 | n2412 ;
  assign n2414 = n232 | n2413 ;
  assign n2415 = n256 | n2414 ;
  assign n2416 = n553 | n2415 ;
  assign n2417 = n339 | n2416 ;
  assign n2418 = n293 | n2417 ;
  assign n2419 = n2128 & n2130 ;
  assign n6024 = ~n2419 ;
  assign n2420 = n2131 & n6024 ;
  assign n6025 = ~n2420 ;
  assign n2422 = n2418 & n6025 ;
  assign n2423 = n552 | n598 ;
  assign n2424 = n332 | n2423 ;
  assign n2425 = n108 | n2424 ;
  assign n2426 = n476 | n2425 ;
  assign n2427 = n293 | n448 ;
  assign n2428 = n996 | n2427 ;
  assign n2429 = n2426 | n2428 ;
  assign n2430 = n2280 | n2429 ;
  assign n2431 = n370 | n2430 ;
  assign n2432 = n2336 | n2431 ;
  assign n2433 = n952 | n2432 ;
  assign n2434 = n356 | n2433 ;
  assign n2435 = n355 | n2434 ;
  assign n2436 = n471 | n2435 ;
  assign n2437 = n221 | n2436 ;
  assign n2438 = n348 | n503 ;
  assign n2439 = n393 | n822 ;
  assign n2440 = n2438 | n2439 ;
  assign n2441 = n2404 | n2440 ;
  assign n6026 = ~n2441 ;
  assign n2442 = n322 & n6026 ;
  assign n6027 = ~n320 ;
  assign n2443 = n6027 & n2442 ;
  assign n6028 = ~n1009 ;
  assign n2444 = n6028 & n2443 ;
  assign n6029 = ~n2437 ;
  assign n2445 = n6029 & n2444 ;
  assign n6030 = ~n162 ;
  assign n2446 = n6030 & n2445 ;
  assign n6031 = ~n325 ;
  assign n2447 = n6031 & n2446 ;
  assign n6032 = ~n212 ;
  assign n2448 = n6032 & n2447 ;
  assign n6033 = ~n255 ;
  assign n2449 = n6033 & n2448 ;
  assign n2450 = n5725 & n2449 ;
  assign n6034 = ~n236 ;
  assign n2451 = n6034 & n2450 ;
  assign n6035 = ~n2125 ;
  assign n2126 = n2123 & n6035 ;
  assign n6036 = ~n2123 ;
  assign n2452 = n6036 & n2125 ;
  assign n2453 = n2126 | n2452 ;
  assign n2454 = n2451 | n2453 ;
  assign n2455 = n2451 & n2453 ;
  assign n2456 = n149 | n1164 ;
  assign n2457 = n225 | n2456 ;
  assign n2458 = n344 | n2457 ;
  assign n2459 = n553 | n2458 ;
  assign n2460 = n173 | n309 ;
  assign n2461 = n367 | n2460 ;
  assign n2462 = n358 | n2461 ;
  assign n2463 = n129 | n2462 ;
  assign n2464 = n2459 | n2463 ;
  assign n2465 = n340 | n2464 ;
  assign n2466 = n457 | n2465 ;
  assign n2467 = n356 | n2466 ;
  assign n2468 = n551 | n2467 ;
  assign n2469 = n151 | n2468 ;
  assign n2470 = n254 | n2427 ;
  assign n2471 = n473 | n2470 ;
  assign n2472 = n2342 | n2471 ;
  assign n2473 = n2469 | n2472 ;
  assign n2474 = n805 | n2473 ;
  assign n2475 = n334 | n2474 ;
  assign n2476 = n206 | n2475 ;
  assign n2477 = n131 | n2476 ;
  assign n2478 = n190 | n2477 ;
  assign n2479 = n120 | n2478 ;
  assign n2480 = n222 | n2479 ;
  assign n2481 = n354 | n2480 ;
  assign n2482 = n444 | n2481 ;
  assign n2483 = n1830 | n2117 ;
  assign n2484 = n2116 | n2483 ;
  assign n2486 = n5980 & n2484 ;
  assign n6037 = ~n2121 ;
  assign n2487 = n6037 & n2486 ;
  assign n6038 = ~n2486 ;
  assign n2488 = n2121 & n6038 ;
  assign n2489 = n2487 | n2488 ;
  assign n6039 = ~n2489 ;
  assign n2490 = n2482 & n6039 ;
  assign n6040 = ~n2482 ;
  assign n2491 = n6040 & n2489 ;
  assign n6041 = ~n2483 ;
  assign n2485 = n2116 & n6041 ;
  assign n6042 = ~n2116 ;
  assign n2492 = n6042 & n2483 ;
  assign n2493 = n2485 | n2492 ;
  assign n2180 = n412 | n625 ;
  assign n2181 = n294 | n2180 ;
  assign n2182 = n353 | n2181 ;
  assign n2185 = n554 | n2184 ;
  assign n2186 = n475 | n2185 ;
  assign n2187 = n1138 | n2186 ;
  assign n2188 = n2182 | n2187 ;
  assign n2189 = n1012 | n2188 ;
  assign n2190 = n769 | n2189 ;
  assign n2191 = n151 | n2190 ;
  assign n2494 = n793 | n1143 ;
  assign n2495 = n940 | n2494 ;
  assign n2496 = n370 | n2495 ;
  assign n2497 = n2399 | n2496 ;
  assign n2498 = n755 | n2497 ;
  assign n2499 = n2191 | n2498 ;
  assign n2500 = n414 | n2499 ;
  assign n2501 = n190 | n2500 ;
  assign n2502 = n355 | n2501 ;
  assign n2503 = n188 | n2502 ;
  assign n2504 = n598 | n2503 ;
  assign n6043 = ~n2504 ;
  assign n2505 = n2493 & n6043 ;
  assign n2506 = n2491 | n2505 ;
  assign n6044 = ~n2490 ;
  assign n2507 = n6044 & n2506 ;
  assign n2509 = n2455 | n2507 ;
  assign n2510 = n2454 & n2509 ;
  assign n6045 = ~n2418 ;
  assign n2421 = n6045 & n2420 ;
  assign n2511 = n2421 | n2422 ;
  assign n2512 = n2510 | n2511 ;
  assign n6046 = ~n2422 ;
  assign n2513 = n6046 & n2512 ;
  assign n6047 = ~n2389 ;
  assign n2391 = n6047 & n2390 ;
  assign n2514 = n2391 | n2392 ;
  assign n2516 = n2513 | n2514 ;
  assign n6048 = ~n2392 ;
  assign n2517 = n6048 & n2516 ;
  assign n2518 = n2361 | n2517 ;
  assign n6049 = ~n2360 ;
  assign n2519 = n6049 & n2518 ;
  assign n2332 = n2330 & n2331 ;
  assign n2520 = n2330 | n2331 ;
  assign n6050 = ~n2332 ;
  assign n2521 = n6050 & n2520 ;
  assign n2523 = n2519 | n2521 ;
  assign n6051 = ~n2333 ;
  assign n2524 = n6051 & n2523 ;
  assign n2525 = n2297 | n2524 ;
  assign n2526 = n2298 & n2525 ;
  assign n6052 = ~n2266 ;
  assign n2268 = n6052 & n2267 ;
  assign n2528 = n2268 | n2269 ;
  assign n2530 = n2526 | n2528 ;
  assign n6053 = ~n2269 ;
  assign n2531 = n6053 & n2530 ;
  assign n2532 = n2230 | n2531 ;
  assign n6054 = ~n2229 ;
  assign n2533 = n6054 & n2532 ;
  assign n2168 = n252 | n326 ;
  assign n2169 = n355 | n2168 ;
  assign n2170 = n323 | n2169 ;
  assign n2171 = n339 | n2170 ;
  assign n2172 = n776 | n2171 ;
  assign n2173 = n224 | n2172 ;
  assign n2174 = n216 | n2173 ;
  assign n2175 = n164 | n2174 ;
  assign n2176 = n204 | n2175 ;
  assign n2177 = n188 | n2176 ;
  assign n2178 = n588 | n2177 ;
  assign n2179 = n752 | n2178 ;
  assign n2198 = n150 | n824 ;
  assign n2199 = n394 | n2198 ;
  assign n2200 = n789 | n2199 ;
  assign n2201 = n2197 | n2200 ;
  assign n2202 = n2191 | n2201 ;
  assign n2203 = n2179 | n2202 ;
  assign n2204 = n2167 | n2203 ;
  assign n2205 = n325 | n2204 ;
  assign n2206 = n226 | n2205 ;
  assign n2207 = n174 | n2206 ;
  assign n2208 = n503 | n2207 ;
  assign n2209 = n364 | n2208 ;
  assign n2210 = n213 | n2209 ;
  assign n732 = n705 & n730 ;
  assign n738 = n732 | n737 ;
  assign n530 = n441 & n528 ;
  assign n544 = n523 & n5689 ;
  assign n6055 = ~n538 ;
  assign n540 = n523 & n6055 ;
  assign n546 = n540 | n545 ;
  assign n6056 = ~n544 ;
  assign n547 = n6056 & n546 ;
  assign n6057 = ~n530 ;
  assign n548 = n6057 & n547 ;
  assign n6058 = ~n547 ;
  assign n549 = n530 & n6058 ;
  assign n550 = n548 | n549 ;
  assign n682 = n674 | n679 ;
  assign n739 = n550 & n682 ;
  assign n6059 = ~n549 ;
  assign n683 = n6059 & n682 ;
  assign n684 = n548 | n683 ;
  assign n740 = n549 | n684 ;
  assign n6060 = ~n739 ;
  assign n741 = n6060 & n740 ;
  assign n742 = n738 & n741 ;
  assign n743 = n738 | n741 ;
  assign n6061 = ~n742 ;
  assign n744 = n6061 & n743 ;
  assign n6062 = ~n924 ;
  assign n926 = n922 & n6062 ;
  assign n6063 = ~n926 ;
  assign n2152 = n6063 & n2151 ;
  assign n2153 = n744 & n2152 ;
  assign n2154 = n744 | n2152 ;
  assign n6064 = ~n2153 ;
  assign n2211 = n6064 & n2154 ;
  assign n6065 = ~n2210 ;
  assign n2212 = n6065 & n2211 ;
  assign n6066 = ~n2211 ;
  assign n2213 = n2210 & n6066 ;
  assign n2534 = n2212 | n2213 ;
  assign n6067 = ~n2534 ;
  assign n2535 = n2533 & n6067 ;
  assign n6068 = ~n2533 ;
  assign n2563 = n6068 & n2534 ;
  assign n2564 = n2535 | n2563 ;
  assign n2565 = n2562 & n2564 ;
  assign n329 = n324 | n328 ;
  assign n330 = n165 | n329 ;
  assign n331 = n323 | n330 ;
  assign n335 = n186 | n334 ;
  assign n336 = n172 | n335 ;
  assign n337 = n333 | n336 ;
  assign n338 = n332 | n337 ;
  assign n343 = n147 | n342 ;
  assign n380 = n346 | n379 ;
  assign n381 = n343 | n380 ;
  assign n382 = n257 | n381 ;
  assign n383 = n341 | n382 ;
  assign n384 = n338 | n383 ;
  assign n385 = n331 | n384 ;
  assign n6069 = ~n385 ;
  assign n386 = n322 & n6069 ;
  assign n387 = n6027 & n386 ;
  assign n388 = n5601 & n387 ;
  assign n389 = n5737 & n388 ;
  assign n6070 = ~n131 ;
  assign n390 = n6070 & n389 ;
  assign n529 = n523 & n528 ;
  assign n531 = n523 | n528 ;
  assign n6071 = ~n529 ;
  assign n532 = n6071 & n531 ;
  assign n6072 = ~n532 ;
  assign n533 = n520 & n6072 ;
  assign n534 = n5510 & n532 ;
  assign n535 = n533 | n534 ;
  assign n6073 = ~n535 ;
  assign n536 = n441 & n6073 ;
  assign n6074 = ~n741 ;
  assign n2155 = n738 & n6074 ;
  assign n6075 = ~n2155 ;
  assign n2156 = n2154 & n6075 ;
  assign n2157 = n684 & n2156 ;
  assign n2158 = n684 | n2156 ;
  assign n6076 = ~n2157 ;
  assign n2159 = n6076 & n2158 ;
  assign n2160 = n536 & n2159 ;
  assign n2161 = n536 | n2159 ;
  assign n6077 = ~n2160 ;
  assign n2162 = n6077 & n2161 ;
  assign n2163 = n390 | n2162 ;
  assign n2164 = n390 & n2162 ;
  assign n6078 = ~n2164 ;
  assign n2165 = n2163 & n6078 ;
  assign n2536 = n2533 | n2534 ;
  assign n6079 = ~n2213 ;
  assign n2537 = n6079 & n2536 ;
  assign n2568 = n2165 | n2537 ;
  assign n2538 = n2164 | n2537 ;
  assign n2539 = n2163 & n2538 ;
  assign n2569 = n6078 & n2539 ;
  assign n6080 = ~n2569 ;
  assign n2570 = n2568 & n6080 ;
  assign n2574 = n5503 & n2560 ;
  assign n6081 = ~n2570 ;
  assign n2575 = n6081 & n2574 ;
  assign n2578 = n2565 | n2575 ;
  assign n6082 = ~n278 ;
  assign n292 = n6082 & n291 ;
  assign n2540 = n405 | n812 ;
  assign n2541 = n186 | n2540 ;
  assign n2542 = n225 | n2541 ;
  assign n2543 = n171 | n2542 ;
  assign n2544 = n365 | n2543 ;
  assign n2545 = n477 | n1138 ;
  assign n2546 = n2342 | n2545 ;
  assign n2547 = n1525 | n2546 ;
  assign n2548 = n2544 | n2547 ;
  assign n2549 = n652 | n2548 ;
  assign n2550 = n146 | n2549 ;
  assign n2551 = n296 | n2550 ;
  assign n2552 = n971 | n2551 ;
  assign n2553 = n551 | n2552 ;
  assign n2554 = n553 | n2553 ;
  assign n2555 = n221 | n2554 ;
  assign n6083 = ~n2555 ;
  assign n2556 = n2539 & n6083 ;
  assign n6084 = ~n2539 ;
  assign n2557 = n6084 & n2555 ;
  assign n2558 = n2556 | n2557 ;
  assign n2579 = n292 & n2558 ;
  assign n2580 = n2578 | n2579 ;
  assign n2581 = n278 & n291 ;
  assign n2231 = n2229 | n2230 ;
  assign n6085 = ~n2531 ;
  assign n2582 = n2231 & n6085 ;
  assign n6086 = ~n2230 ;
  assign n2583 = n6086 & n2533 ;
  assign n2584 = n2582 | n2583 ;
  assign n6087 = ~n2528 ;
  assign n2529 = n2526 & n6087 ;
  assign n6088 = ~n2526 ;
  assign n2588 = n6088 & n2528 ;
  assign n2589 = n2529 | n2588 ;
  assign n2591 = n2584 & n2589 ;
  assign n6089 = ~n2297 ;
  assign n2527 = n6089 & n2526 ;
  assign n2299 = n6089 & n2298 ;
  assign n2593 = n2299 | n2524 ;
  assign n6090 = ~n2527 ;
  assign n2594 = n6090 & n2593 ;
  assign n6091 = ~n2594 ;
  assign n2595 = n2589 & n6091 ;
  assign n6092 = ~n2519 ;
  assign n2522 = n6092 & n2521 ;
  assign n6093 = ~n2521 ;
  assign n2597 = n2519 & n6093 ;
  assign n2598 = n2522 | n2597 ;
  assign n2600 = n6091 & n2598 ;
  assign n2362 = n2360 | n2361 ;
  assign n6094 = ~n2517 ;
  assign n2603 = n2362 & n6094 ;
  assign n6095 = ~n2361 ;
  assign n2604 = n6095 & n2519 ;
  assign n2605 = n2603 | n2604 ;
  assign n2606 = n2598 & n2605 ;
  assign n6096 = ~n2514 ;
  assign n2515 = n2513 & n6096 ;
  assign n6097 = ~n2513 ;
  assign n2610 = n6097 & n2514 ;
  assign n2611 = n2515 | n2610 ;
  assign n2613 = n2605 & n2611 ;
  assign n2615 = n2510 & n2511 ;
  assign n6098 = ~n2615 ;
  assign n2616 = n2512 & n6098 ;
  assign n2619 = n2611 & n2616 ;
  assign n6099 = ~n2455 ;
  assign n2621 = n2454 & n6099 ;
  assign n2622 = n2507 | n2621 ;
  assign n2623 = n6099 & n2510 ;
  assign n6100 = ~n2623 ;
  assign n2624 = n2622 & n6100 ;
  assign n6101 = ~n2624 ;
  assign n2625 = n2616 & n6101 ;
  assign n6102 = ~n2491 ;
  assign n2508 = n6102 & n2507 ;
  assign n2620 = n2490 | n2491 ;
  assign n6103 = ~n2505 ;
  assign n2629 = n6103 & n2620 ;
  assign n2630 = n2508 | n2629 ;
  assign n6104 = ~n2493 ;
  assign n2632 = n6104 & n2504 ;
  assign n2633 = n2505 | n2632 ;
  assign n6105 = ~n2633 ;
  assign n2634 = n2624 & n6105 ;
  assign n6106 = ~n2634 ;
  assign n2635 = n2630 & n6106 ;
  assign n6107 = ~n2616 ;
  assign n2636 = n6107 & n2624 ;
  assign n6108 = ~n2636 ;
  assign n2637 = n2635 & n6108 ;
  assign n2638 = n2625 | n2637 ;
  assign n2639 = n2611 | n2616 ;
  assign n2640 = n2638 & n2639 ;
  assign n2642 = n2619 | n2640 ;
  assign n6109 = ~n2605 ;
  assign n2612 = n6109 & n2611 ;
  assign n6110 = ~n2611 ;
  assign n2644 = n2605 & n6110 ;
  assign n2645 = n2612 | n2644 ;
  assign n2647 = n2642 & n2645 ;
  assign n2648 = n2613 | n2647 ;
  assign n2608 = n2598 | n2605 ;
  assign n6111 = ~n2606 ;
  assign n2649 = n6111 & n2608 ;
  assign n2651 = n2648 & n2649 ;
  assign n2652 = n2606 | n2651 ;
  assign n6112 = ~n2598 ;
  assign n2602 = n2594 & n6112 ;
  assign n2653 = n2600 | n2602 ;
  assign n6113 = ~n2653 ;
  assign n2655 = n2652 & n6113 ;
  assign n2656 = n2600 | n2655 ;
  assign n6114 = ~n2589 ;
  assign n2596 = n6114 & n2594 ;
  assign n2657 = n2595 | n2596 ;
  assign n6115 = ~n2657 ;
  assign n2659 = n2656 & n6115 ;
  assign n2660 = n2595 | n2659 ;
  assign n2592 = n2584 | n2589 ;
  assign n6116 = ~n2591 ;
  assign n2661 = n6116 & n2592 ;
  assign n2663 = n2660 & n2661 ;
  assign n2664 = n2591 | n2663 ;
  assign n6117 = ~n2584 ;
  assign n2587 = n2564 & n6117 ;
  assign n6118 = ~n2564 ;
  assign n2665 = n6118 & n2584 ;
  assign n2666 = n2587 | n2665 ;
  assign n2668 = n2664 & n2666 ;
  assign n2669 = n2564 & n2584 ;
  assign n2670 = n2668 | n2669 ;
  assign n2572 = n2564 & n2570 ;
  assign n2671 = n2564 | n2570 ;
  assign n6119 = ~n2572 ;
  assign n2672 = n6119 & n2671 ;
  assign n6120 = ~n2672 ;
  assign n2673 = n2670 & n6120 ;
  assign n2674 = n2564 & n6081 ;
  assign n2675 = n2673 | n2674 ;
  assign n6121 = ~n2558 ;
  assign n2573 = n6121 & n2570 ;
  assign n2676 = n2558 & n6081 ;
  assign n2677 = n2573 | n2676 ;
  assign n6122 = ~n2677 ;
  assign n2678 = n2675 & n6122 ;
  assign n6123 = ~n2675 ;
  assign n2679 = n6123 & n2677 ;
  assign n2680 = n2678 | n2679 ;
  assign n6124 = ~n2680 ;
  assign n2681 = n2581 & n6124 ;
  assign n2682 = n2580 | n2681 ;
  assign n6125 = ~n2682 ;
  assign n2683 = n274 & n6125 ;
  assign n2684 = n5721 & n2682 ;
  assign n2685 = n2683 | n2684 ;
  assign n681 = n672 & n5550 ;
  assign n2686 = n5514 & n677 ;
  assign n2687 = n681 | n2686 ;
  assign n2688 = n2633 & n2687 ;
  assign n6126 = ~n2688 ;
  assign n2689 = n523 & n6126 ;
  assign n680 = n528 | n677 ;
  assign n2691 = n528 & n677 ;
  assign n6127 = ~n2691 ;
  assign n2692 = n680 & n6127 ;
  assign n6128 = ~n2687 ;
  assign n2693 = n6128 & n2692 ;
  assign n2707 = n2633 & n2693 ;
  assign n2699 = n6072 & n2687 ;
  assign n2708 = n2630 & n2699 ;
  assign n2709 = n2707 | n2708 ;
  assign n2690 = n2630 | n2633 ;
  assign n2710 = n2630 & n2633 ;
  assign n6129 = ~n2710 ;
  assign n2711 = n2690 & n6129 ;
  assign n2713 = n532 & n2687 ;
  assign n2715 = n2711 & n2713 ;
  assign n2716 = n2709 | n2715 ;
  assign n6130 = ~n2716 ;
  assign n2717 = n523 & n6130 ;
  assign n2718 = n5542 & n2716 ;
  assign n2719 = n2717 | n2718 ;
  assign n6131 = ~n2719 ;
  assign n2720 = n2689 & n6131 ;
  assign n6132 = ~n2689 ;
  assign n2721 = n6132 & n2719 ;
  assign n2722 = n2720 | n2721 ;
  assign n866 = n851 & n5512 ;
  assign n2730 = n5554 & n859 ;
  assign n2731 = n866 | n2730 ;
  assign n1058 = n851 | n1052 ;
  assign n2723 = n851 & n1052 ;
  assign n6133 = ~n2723 ;
  assign n2724 = n1058 & n6133 ;
  assign n865 = n672 | n859 ;
  assign n2725 = n672 & n859 ;
  assign n6134 = ~n2725 ;
  assign n2726 = n865 & n6134 ;
  assign n6135 = ~n2724 ;
  assign n2732 = n6135 & n2726 ;
  assign n6136 = ~n2731 ;
  assign n2733 = n6136 & n2732 ;
  assign n2735 = n6101 & n2733 ;
  assign n2742 = n6135 & n2731 ;
  assign n2755 = n2616 & n2742 ;
  assign n6137 = ~n2726 ;
  assign n2748 = n2724 & n6137 ;
  assign n2756 = n2611 & n2748 ;
  assign n2757 = n2755 | n2756 ;
  assign n2758 = n2735 | n2757 ;
  assign n2727 = n2724 & n2726 ;
  assign n6138 = ~n2642 ;
  assign n2643 = n2639 & n6138 ;
  assign n6139 = ~n2619 ;
  assign n2641 = n6139 & n2639 ;
  assign n6140 = ~n2641 ;
  assign n2759 = n2638 & n6140 ;
  assign n2760 = n2643 | n2759 ;
  assign n2761 = n2727 & n2760 ;
  assign n2762 = n2758 | n2761 ;
  assign n2763 = n672 & n2762 ;
  assign n2764 = n672 | n2762 ;
  assign n6141 = ~n2763 ;
  assign n2765 = n6141 & n2764 ;
  assign n2766 = n2722 & n2765 ;
  assign n2767 = n2633 & n2724 ;
  assign n6142 = ~n2767 ;
  assign n2768 = n672 & n6142 ;
  assign n2728 = n2711 & n2727 ;
  assign n2769 = n2633 & n2742 ;
  assign n2770 = n2630 & n2748 ;
  assign n2771 = n2769 | n2770 ;
  assign n2772 = n2728 | n2771 ;
  assign n6143 = ~n2772 ;
  assign n2773 = n672 & n6143 ;
  assign n2774 = n5514 & n2772 ;
  assign n2775 = n2773 | n2774 ;
  assign n2776 = n2768 & n2775 ;
  assign n2751 = n6101 & n2748 ;
  assign n2777 = n2633 & n2733 ;
  assign n2778 = n2630 & n2742 ;
  assign n2779 = n2777 | n2778 ;
  assign n2780 = n2751 | n2779 ;
  assign n2781 = n2630 & n6105 ;
  assign n2782 = n6101 & n2781 ;
  assign n6144 = ~n2781 ;
  assign n2783 = n2624 & n6144 ;
  assign n2784 = n2782 | n2783 ;
  assign n6145 = ~n2784 ;
  assign n2785 = n2727 & n6145 ;
  assign n2786 = n2780 | n2785 ;
  assign n2787 = n672 & n2786 ;
  assign n2788 = n672 | n2786 ;
  assign n6146 = ~n2787 ;
  assign n2789 = n6146 & n2788 ;
  assign n2790 = n2776 & n2789 ;
  assign n2792 = n2688 & n2790 ;
  assign n2791 = n6126 & n2790 ;
  assign n6147 = ~n2790 ;
  assign n2793 = n2688 & n6147 ;
  assign n2794 = n2791 | n2793 ;
  assign n2736 = n2630 & n2733 ;
  assign n2752 = n2616 & n2748 ;
  assign n2795 = n2736 | n2752 ;
  assign n2796 = n6101 & n2742 ;
  assign n2797 = n2795 | n2796 ;
  assign n2798 = n2625 | n2636 ;
  assign n2799 = n2635 & n2798 ;
  assign n2800 = n2636 | n2638 ;
  assign n6148 = ~n2799 ;
  assign n2801 = n6148 & n2800 ;
  assign n6149 = ~n2801 ;
  assign n2802 = n2727 & n6149 ;
  assign n2805 = n2797 | n2802 ;
  assign n6150 = ~n2805 ;
  assign n2806 = n672 & n6150 ;
  assign n2807 = n5514 & n2805 ;
  assign n2808 = n2806 | n2807 ;
  assign n2810 = n2794 & n2808 ;
  assign n2811 = n2792 | n2810 ;
  assign n2812 = n2722 | n2765 ;
  assign n6151 = ~n2766 ;
  assign n2813 = n6151 & n2812 ;
  assign n2815 = n2811 & n2813 ;
  assign n2816 = n2766 | n2815 ;
  assign n2739 = n2616 & n2733 ;
  assign n2743 = n2611 & n2742 ;
  assign n2817 = n2739 | n2743 ;
  assign n2818 = n2605 & n2748 ;
  assign n2819 = n2817 | n2818 ;
  assign n2646 = n6138 & n2645 ;
  assign n6152 = ~n2645 ;
  assign n2820 = n2642 & n6152 ;
  assign n2821 = n2646 | n2820 ;
  assign n2822 = n2727 & n2821 ;
  assign n2825 = n2819 | n2822 ;
  assign n6153 = ~n2825 ;
  assign n2826 = n672 & n6153 ;
  assign n2827 = n5514 & n2825 ;
  assign n2828 = n2826 | n2827 ;
  assign n2829 = n2689 & n2719 ;
  assign n2700 = n6101 & n2699 ;
  assign n2838 = n2630 & n2693 ;
  assign n2830 = n532 & n6128 ;
  assign n6154 = ~n2692 ;
  assign n2831 = n6154 & n2830 ;
  assign n2839 = n2633 & n2831 ;
  assign n2840 = n2838 | n2839 ;
  assign n2841 = n2700 | n2840 ;
  assign n2842 = n2713 & n6145 ;
  assign n2843 = n2841 | n2842 ;
  assign n2844 = n523 & n2843 ;
  assign n2845 = n523 | n2843 ;
  assign n6155 = ~n2844 ;
  assign n2846 = n6155 & n2845 ;
  assign n2847 = n2829 & n2846 ;
  assign n2848 = n2829 | n2846 ;
  assign n6156 = ~n2847 ;
  assign n2849 = n6156 & n2848 ;
  assign n2850 = n2828 & n2849 ;
  assign n2851 = n2828 | n2849 ;
  assign n6157 = ~n2850 ;
  assign n2852 = n6157 & n2851 ;
  assign n6158 = ~n2816 ;
  assign n2853 = n6158 & n2852 ;
  assign n6159 = ~n2852 ;
  assign n2854 = n2816 & n6159 ;
  assign n2855 = n2853 | n2854 ;
  assign n1057 = n1043 & n5595 ;
  assign n2856 = n5647 & n1052 ;
  assign n2857 = n1057 | n2856 ;
  assign n1238 = n274 & n5722 ;
  assign n2858 = n5721 & n1229 ;
  assign n2859 = n1238 | n2858 ;
  assign n6160 = ~n2857 ;
  assign n2860 = n6160 & n2859 ;
  assign n2861 = n2589 & n2860 ;
  assign n1237 = n1043 | n1229 ;
  assign n2867 = n1043 & n1229 ;
  assign n6161 = ~n2867 ;
  assign n2868 = n1237 & n6161 ;
  assign n6162 = ~n2859 ;
  assign n2869 = n2857 & n6162 ;
  assign n6163 = ~n2868 ;
  assign n2870 = n6163 & n2869 ;
  assign n2885 = n2598 & n2870 ;
  assign n2879 = n6162 & n2868 ;
  assign n2886 = n6091 & n2879 ;
  assign n2887 = n2885 | n2886 ;
  assign n2888 = n2861 | n2887 ;
  assign n2658 = n2656 | n2657 ;
  assign n2889 = n2656 & n2657 ;
  assign n6164 = ~n2889 ;
  assign n2890 = n2658 & n6164 ;
  assign n2891 = n2857 & n2859 ;
  assign n6165 = ~n2890 ;
  assign n2896 = n6165 & n2891 ;
  assign n2897 = n2888 | n2896 ;
  assign n2898 = n1052 & n2897 ;
  assign n2899 = n1052 | n2897 ;
  assign n6166 = ~n2898 ;
  assign n2900 = n6166 & n2899 ;
  assign n2902 = n2855 & n2900 ;
  assign n2871 = n2605 & n2870 ;
  assign n2880 = n2598 & n2879 ;
  assign n2903 = n2871 | n2880 ;
  assign n2904 = n6091 & n2860 ;
  assign n2905 = n2903 | n2904 ;
  assign n2654 = n2652 | n2653 ;
  assign n2906 = n2652 & n2653 ;
  assign n6167 = ~n2906 ;
  assign n2907 = n2654 & n6167 ;
  assign n6168 = ~n2907 ;
  assign n2908 = n2891 & n6168 ;
  assign n2912 = n2905 | n2908 ;
  assign n6169 = ~n2912 ;
  assign n2913 = n1052 & n6169 ;
  assign n2914 = n5595 & n2912 ;
  assign n2915 = n2913 | n2914 ;
  assign n6170 = ~n2811 ;
  assign n2814 = n6170 & n2813 ;
  assign n6171 = ~n2813 ;
  assign n2916 = n2811 & n6171 ;
  assign n2917 = n2814 | n2916 ;
  assign n2919 = n2915 & n2917 ;
  assign n6172 = ~n2794 ;
  assign n2809 = n6172 & n2808 ;
  assign n6173 = ~n2808 ;
  assign n2920 = n2794 & n6173 ;
  assign n2921 = n2809 | n2920 ;
  assign n2863 = n2598 & n2860 ;
  assign n2922 = n2611 & n2870 ;
  assign n2923 = n2605 & n2879 ;
  assign n2924 = n2922 | n2923 ;
  assign n2925 = n2863 | n2924 ;
  assign n6174 = ~n2648 ;
  assign n2650 = n6174 & n2649 ;
  assign n6175 = ~n2649 ;
  assign n2926 = n2648 & n6175 ;
  assign n2927 = n2650 | n2926 ;
  assign n2928 = n2891 & n2927 ;
  assign n2929 = n2925 | n2928 ;
  assign n2930 = n1052 & n2929 ;
  assign n2931 = n1052 | n2929 ;
  assign n6176 = ~n2930 ;
  assign n2932 = n6176 & n2931 ;
  assign n2934 = n2921 & n2932 ;
  assign n2895 = n2821 & n2891 ;
  assign n2873 = n2616 & n2870 ;
  assign n2882 = n2611 & n2879 ;
  assign n2935 = n2873 | n2882 ;
  assign n2936 = n2605 & n2860 ;
  assign n2937 = n2935 | n2936 ;
  assign n2938 = n2895 | n2937 ;
  assign n6177 = ~n2938 ;
  assign n2939 = n1052 & n6177 ;
  assign n2940 = n5595 & n2938 ;
  assign n2941 = n2939 | n2940 ;
  assign n2942 = n2776 | n2789 ;
  assign n2943 = n6147 & n2942 ;
  assign n2945 = n2941 & n2943 ;
  assign n2946 = n2768 | n2775 ;
  assign n6178 = ~n2776 ;
  assign n2947 = n6178 & n2946 ;
  assign n2874 = n6101 & n2870 ;
  assign n2948 = n2611 & n2860 ;
  assign n2949 = n2616 & n2879 ;
  assign n2950 = n2948 | n2949 ;
  assign n2951 = n2874 | n2950 ;
  assign n2952 = n2760 & n2891 ;
  assign n2953 = n2951 | n2952 ;
  assign n2954 = n1052 & n2953 ;
  assign n2955 = n1052 | n2953 ;
  assign n6179 = ~n2954 ;
  assign n2956 = n6179 & n2955 ;
  assign n2957 = n2947 & n2956 ;
  assign n2894 = n2711 & n2891 ;
  assign n2958 = n2630 & n2860 ;
  assign n2959 = n2633 & n2879 ;
  assign n2960 = n2958 | n2959 ;
  assign n2961 = n2894 | n2960 ;
  assign n6180 = ~n2961 ;
  assign n2962 = n1052 & n6180 ;
  assign n2963 = n5595 & n2961 ;
  assign n2964 = n2962 | n2963 ;
  assign n2965 = n2633 & n2859 ;
  assign n6181 = ~n2965 ;
  assign n2966 = n1052 & n6181 ;
  assign n2968 = n2964 & n2966 ;
  assign n2865 = n6101 & n2860 ;
  assign n2969 = n2633 & n2870 ;
  assign n2970 = n2630 & n2879 ;
  assign n2971 = n2969 | n2970 ;
  assign n2972 = n2865 | n2971 ;
  assign n2973 = n6145 & n2891 ;
  assign n2974 = n2972 | n2973 ;
  assign n2975 = n1052 & n2974 ;
  assign n2976 = n1052 | n2974 ;
  assign n6182 = ~n2975 ;
  assign n2977 = n6182 & n2976 ;
  assign n2978 = n2968 & n2977 ;
  assign n2980 = n2767 & n2978 ;
  assign n2979 = n6142 & n2978 ;
  assign n6183 = ~n2978 ;
  assign n2981 = n2767 & n6183 ;
  assign n2982 = n2979 | n2981 ;
  assign n2893 = n6149 & n2891 ;
  assign n2862 = n2616 & n2860 ;
  assign n2872 = n2630 & n2870 ;
  assign n2983 = n2862 | n2872 ;
  assign n2984 = n6101 & n2879 ;
  assign n2985 = n2983 | n2984 ;
  assign n2986 = n2893 | n2985 ;
  assign n6184 = ~n2986 ;
  assign n2987 = n1052 & n6184 ;
  assign n2988 = n5595 & n2986 ;
  assign n2989 = n2987 | n2988 ;
  assign n2991 = n2982 & n2989 ;
  assign n2992 = n2980 | n2991 ;
  assign n2993 = n2947 | n2956 ;
  assign n6185 = ~n2957 ;
  assign n2994 = n6185 & n2993 ;
  assign n2996 = n2992 & n2994 ;
  assign n2997 = n2957 | n2996 ;
  assign n6186 = ~n2941 ;
  assign n2944 = n6186 & n2943 ;
  assign n6187 = ~n2943 ;
  assign n2998 = n2941 & n6187 ;
  assign n2999 = n2944 | n2998 ;
  assign n3001 = n2997 & n2999 ;
  assign n3002 = n2945 | n3001 ;
  assign n6188 = ~n2921 ;
  assign n2933 = n6188 & n2932 ;
  assign n6189 = ~n2932 ;
  assign n3003 = n2921 & n6189 ;
  assign n3004 = n2933 | n3003 ;
  assign n3006 = n3002 & n3004 ;
  assign n3007 = n2934 | n3006 ;
  assign n6190 = ~n2915 ;
  assign n2918 = n6190 & n2917 ;
  assign n6191 = ~n2917 ;
  assign n3008 = n2915 & n6191 ;
  assign n3009 = n2918 | n3008 ;
  assign n3011 = n3007 & n3009 ;
  assign n3012 = n2919 | n3011 ;
  assign n6192 = ~n2855 ;
  assign n2901 = n6192 & n2900 ;
  assign n6193 = ~n2900 ;
  assign n3013 = n2855 & n6193 ;
  assign n3014 = n2901 | n3013 ;
  assign n3016 = n3012 & n3014 ;
  assign n3017 = n2902 | n3016 ;
  assign n2740 = n2611 & n2733 ;
  assign n2744 = n2605 & n2742 ;
  assign n3018 = n2740 | n2744 ;
  assign n3019 = n2598 & n2748 ;
  assign n3020 = n3018 | n3019 ;
  assign n3021 = n2727 & n2927 ;
  assign n3022 = n3020 | n3021 ;
  assign n6194 = ~n3022 ;
  assign n3023 = n672 & n6194 ;
  assign n3024 = n5514 & n3022 ;
  assign n3025 = n3023 | n3024 ;
  assign n2804 = n2713 & n6149 ;
  assign n2701 = n2616 & n2699 ;
  assign n2832 = n2630 & n2831 ;
  assign n3026 = n2701 | n2832 ;
  assign n3027 = n6101 & n2693 ;
  assign n3028 = n3026 | n3027 ;
  assign n3029 = n2804 | n3028 ;
  assign n6195 = ~n3029 ;
  assign n3030 = n523 & n6195 ;
  assign n3031 = n5542 & n3029 ;
  assign n3032 = n3030 | n3031 ;
  assign n3033 = n523 & n2633 ;
  assign n3034 = n2847 | n3033 ;
  assign n3035 = n2847 & n3033 ;
  assign n6196 = ~n3035 ;
  assign n3036 = n3034 & n6196 ;
  assign n6197 = ~n3036 ;
  assign n3037 = n3032 & n6197 ;
  assign n3038 = n3032 & n3034 ;
  assign n3039 = n3035 | n3038 ;
  assign n6198 = ~n3039 ;
  assign n3040 = n3034 & n6198 ;
  assign n3041 = n3037 | n3040 ;
  assign n6199 = ~n3041 ;
  assign n3042 = n3025 & n6199 ;
  assign n6200 = ~n3025 ;
  assign n3043 = n6200 & n3041 ;
  assign n3044 = n3042 | n3043 ;
  assign n3045 = n2816 & n2852 ;
  assign n3046 = n2850 | n3045 ;
  assign n3047 = n3044 | n3046 ;
  assign n3048 = n3044 & n3046 ;
  assign n6201 = ~n3048 ;
  assign n3049 = n3047 & n6201 ;
  assign n2864 = n2584 & n2860 ;
  assign n3052 = n6091 & n2870 ;
  assign n3053 = n2589 & n2879 ;
  assign n3054 = n3052 | n3053 ;
  assign n3055 = n2864 | n3054 ;
  assign n6202 = ~n2660 ;
  assign n2662 = n6202 & n2661 ;
  assign n6203 = ~n2661 ;
  assign n3050 = n2660 & n6203 ;
  assign n3051 = n2662 | n3050 ;
  assign n3056 = n2891 & n3051 ;
  assign n3057 = n3055 | n3056 ;
  assign n3058 = n1052 & n3057 ;
  assign n3059 = n1052 | n3057 ;
  assign n6204 = ~n3058 ;
  assign n3060 = n6204 & n3059 ;
  assign n6205 = ~n3049 ;
  assign n3061 = n6205 & n3060 ;
  assign n6206 = ~n3060 ;
  assign n3063 = n3049 & n6206 ;
  assign n3064 = n3061 | n3063 ;
  assign n6207 = ~n3064 ;
  assign n3065 = n3017 & n6207 ;
  assign n6208 = ~n3017 ;
  assign n3066 = n6208 & n3064 ;
  assign n3067 = n3065 | n3066 ;
  assign n3068 = n2685 | n3067 ;
  assign n3069 = n2685 & n3067 ;
  assign n6209 = ~n3069 ;
  assign n3070 = n3068 & n6209 ;
  assign n6210 = ~n3014 ;
  assign n3015 = n3012 & n6210 ;
  assign n6211 = ~n3012 ;
  assign n3071 = n6211 & n3014 ;
  assign n3072 = n3015 | n3071 ;
  assign n2576 = n2564 & n2574 ;
  assign n2586 = n2562 & n2584 ;
  assign n3073 = n2576 | n2586 ;
  assign n3074 = n292 & n6081 ;
  assign n3075 = n3073 | n3074 ;
  assign n6212 = ~n2670 ;
  assign n3076 = n6212 & n2672 ;
  assign n3077 = n2673 | n3076 ;
  assign n6213 = ~n3077 ;
  assign n3078 = n2581 & n6213 ;
  assign n3080 = n3075 | n3078 ;
  assign n6214 = ~n3080 ;
  assign n3081 = n274 & n6214 ;
  assign n3082 = n5721 & n3080 ;
  assign n3083 = n3081 | n3082 ;
  assign n3084 = n3072 & n3083 ;
  assign n3085 = n3072 | n3083 ;
  assign n6215 = ~n3084 ;
  assign n3086 = n6215 & n3085 ;
  assign n3010 = n3007 | n3009 ;
  assign n6216 = ~n3011 ;
  assign n3087 = n3010 & n6216 ;
  assign n2566 = n292 & n2564 ;
  assign n3088 = n2574 & n2584 ;
  assign n3089 = n2562 & n2589 ;
  assign n3090 = n3088 | n3089 ;
  assign n3091 = n2566 | n3090 ;
  assign n6217 = ~n2664 ;
  assign n2667 = n6217 & n2666 ;
  assign n6218 = ~n2666 ;
  assign n3092 = n2664 & n6218 ;
  assign n3093 = n2667 | n3092 ;
  assign n3094 = n2581 & n3093 ;
  assign n3095 = n3091 | n3094 ;
  assign n3096 = n274 & n3095 ;
  assign n3097 = n274 | n3095 ;
  assign n6219 = ~n3096 ;
  assign n3098 = n6219 & n3097 ;
  assign n3100 = n3087 & n3098 ;
  assign n6220 = ~n3004 ;
  assign n3005 = n3002 & n6220 ;
  assign n6221 = ~n3002 ;
  assign n3101 = n6221 & n3004 ;
  assign n3102 = n3005 | n3101 ;
  assign n2585 = n292 & n2584 ;
  assign n3103 = n2574 & n2589 ;
  assign n3104 = n2562 & n6091 ;
  assign n3105 = n3103 | n3104 ;
  assign n3106 = n2585 | n3105 ;
  assign n3107 = n2581 & n3051 ;
  assign n3108 = n3106 | n3107 ;
  assign n3109 = n274 & n3108 ;
  assign n3110 = n274 | n3108 ;
  assign n6222 = ~n3109 ;
  assign n3111 = n6222 & n3110 ;
  assign n3113 = n3102 & n3111 ;
  assign n3000 = n2997 | n2999 ;
  assign n6223 = ~n3001 ;
  assign n3114 = n3000 & n6223 ;
  assign n2590 = n292 & n2589 ;
  assign n3115 = n2574 & n6091 ;
  assign n3116 = n2562 & n2598 ;
  assign n3117 = n3115 | n3116 ;
  assign n3118 = n2590 | n3117 ;
  assign n3119 = n2581 & n6165 ;
  assign n3120 = n3118 | n3119 ;
  assign n3121 = n274 & n3120 ;
  assign n3122 = n274 | n3120 ;
  assign n6224 = ~n3121 ;
  assign n3123 = n6224 & n3122 ;
  assign n3125 = n3114 & n3123 ;
  assign n2910 = n2581 & n6168 ;
  assign n2601 = n2574 & n2598 ;
  assign n2607 = n2562 & n2605 ;
  assign n3126 = n2601 | n2607 ;
  assign n3127 = n292 & n6091 ;
  assign n3128 = n3126 | n3127 ;
  assign n3129 = n2910 | n3128 ;
  assign n6225 = ~n3129 ;
  assign n3130 = n274 & n6225 ;
  assign n3131 = n5721 & n3129 ;
  assign n3132 = n3130 | n3131 ;
  assign n6226 = ~n2992 ;
  assign n2995 = n6226 & n2994 ;
  assign n6227 = ~n2994 ;
  assign n3133 = n2992 & n6227 ;
  assign n3134 = n2995 | n3133 ;
  assign n3135 = n3132 & n3134 ;
  assign n2990 = n2982 | n2989 ;
  assign n6228 = ~n2991 ;
  assign n3136 = n2990 & n6228 ;
  assign n2599 = n292 & n2598 ;
  assign n3137 = n2574 & n2605 ;
  assign n3138 = n2562 & n2611 ;
  assign n3139 = n3137 | n3138 ;
  assign n3140 = n2599 | n3139 ;
  assign n3141 = n2581 & n2927 ;
  assign n3142 = n3140 | n3141 ;
  assign n3143 = n274 & n3142 ;
  assign n3144 = n274 | n3142 ;
  assign n6229 = ~n3143 ;
  assign n3145 = n6229 & n3144 ;
  assign n3147 = n3136 & n3145 ;
  assign n2823 = n2581 & n2821 ;
  assign n2614 = n2574 & n2611 ;
  assign n2618 = n2562 & n2616 ;
  assign n3148 = n2614 | n2618 ;
  assign n3149 = n292 & n2605 ;
  assign n3150 = n3148 | n3149 ;
  assign n3151 = n2823 | n3150 ;
  assign n6230 = ~n3151 ;
  assign n3152 = n274 & n6230 ;
  assign n3153 = n5721 & n3151 ;
  assign n3154 = n3152 | n3153 ;
  assign n3155 = n2968 | n2977 ;
  assign n3156 = n6183 & n3155 ;
  assign n3157 = n3154 & n3156 ;
  assign n6231 = ~n2964 ;
  assign n2967 = n6231 & n2966 ;
  assign n6232 = ~n2966 ;
  assign n3158 = n2964 & n6232 ;
  assign n3159 = n2967 | n3158 ;
  assign n2628 = n2562 & n6101 ;
  assign n3160 = n292 & n2611 ;
  assign n3161 = n2574 & n2616 ;
  assign n3162 = n3160 | n3161 ;
  assign n3163 = n2628 | n3162 ;
  assign n3164 = n2581 & n2760 ;
  assign n3165 = n3163 | n3164 ;
  assign n3166 = n274 & n3165 ;
  assign n3167 = n274 | n3165 ;
  assign n6233 = ~n3166 ;
  assign n3168 = n6233 & n3167 ;
  assign n3169 = n3159 & n3168 ;
  assign n3170 = n291 & n2633 ;
  assign n6234 = ~n3170 ;
  assign n3171 = n274 & n6234 ;
  assign n2712 = n2581 & n2711 ;
  assign n3172 = n292 & n2630 ;
  assign n3173 = n2574 & n2633 ;
  assign n3174 = n3172 | n3173 ;
  assign n3175 = n2712 | n3174 ;
  assign n6235 = ~n3175 ;
  assign n3176 = n274 & n6235 ;
  assign n3177 = n5721 & n3175 ;
  assign n3178 = n3176 | n3177 ;
  assign n3179 = n3171 & n3178 ;
  assign n2627 = n292 & n6101 ;
  assign n3180 = n2574 & n2630 ;
  assign n3181 = n2562 & n2633 ;
  assign n3182 = n3180 | n3181 ;
  assign n3183 = n2627 | n3182 ;
  assign n3184 = n2581 & n6145 ;
  assign n3185 = n3183 | n3184 ;
  assign n3186 = n274 & n3185 ;
  assign n3187 = n274 | n3185 ;
  assign n6236 = ~n3186 ;
  assign n3188 = n6236 & n3187 ;
  assign n3189 = n3179 & n3188 ;
  assign n3190 = n2965 & n3189 ;
  assign n3191 = n2965 | n3189 ;
  assign n6237 = ~n3190 ;
  assign n3192 = n6237 & n3191 ;
  assign n2803 = n2581 & n6149 ;
  assign n2617 = n292 & n2616 ;
  assign n2631 = n2562 & n2630 ;
  assign n3193 = n2617 | n2631 ;
  assign n3194 = n2574 & n6101 ;
  assign n3195 = n3193 | n3194 ;
  assign n3196 = n2803 | n3195 ;
  assign n6238 = ~n3196 ;
  assign n3197 = n274 & n6238 ;
  assign n3198 = n5721 & n3196 ;
  assign n3199 = n3197 | n3198 ;
  assign n3201 = n3192 & n3199 ;
  assign n3202 = n3190 | n3201 ;
  assign n3203 = n3159 | n3168 ;
  assign n6239 = ~n3169 ;
  assign n3204 = n6239 & n3203 ;
  assign n3205 = n3202 & n3204 ;
  assign n3206 = n3169 | n3205 ;
  assign n3207 = n3154 | n3156 ;
  assign n6240 = ~n3157 ;
  assign n3208 = n6240 & n3207 ;
  assign n3210 = n3206 & n3208 ;
  assign n3211 = n3157 | n3210 ;
  assign n3146 = n3136 | n3145 ;
  assign n6241 = ~n3147 ;
  assign n3212 = n3146 & n6241 ;
  assign n3214 = n3211 & n3212 ;
  assign n3215 = n3147 | n3214 ;
  assign n3216 = n3132 | n3134 ;
  assign n6242 = ~n3135 ;
  assign n3217 = n6242 & n3216 ;
  assign n3219 = n3215 & n3217 ;
  assign n3220 = n3135 | n3219 ;
  assign n6243 = ~n3114 ;
  assign n3124 = n6243 & n3123 ;
  assign n6244 = ~n3123 ;
  assign n3221 = n3114 & n6244 ;
  assign n3222 = n3124 | n3221 ;
  assign n3224 = n3220 & n3222 ;
  assign n3225 = n3125 | n3224 ;
  assign n6245 = ~n3102 ;
  assign n3112 = n6245 & n3111 ;
  assign n6246 = ~n3111 ;
  assign n3226 = n3102 & n6246 ;
  assign n3227 = n3112 | n3226 ;
  assign n3229 = n3225 & n3227 ;
  assign n3230 = n3113 | n3229 ;
  assign n6247 = ~n3087 ;
  assign n3099 = n6247 & n3098 ;
  assign n6248 = ~n3098 ;
  assign n3231 = n3087 & n6248 ;
  assign n3232 = n3099 | n3231 ;
  assign n3233 = n3230 & n3232 ;
  assign n3234 = n3100 | n3233 ;
  assign n3236 = n3086 & n3234 ;
  assign n3237 = n3084 | n3236 ;
  assign n6249 = ~n3237 ;
  assign n3238 = n3070 & n6249 ;
  assign n6250 = ~n3070 ;
  assign n3239 = n6250 & n3237 ;
  assign n3240 = n3238 | n3239 ;
  assign n3241 = x[0] & n5473 ;
  assign n6251 = ~n3241 ;
  assign n3242 = x[1] & n6251 ;
  assign n6252 = ~x[1] ;
  assign n3243 = n6252 & n3241 ;
  assign n3244 = n3242 | n3243 ;
  assign n3245 = n287 | n3244 ;
  assign n3246 = n287 & n3244 ;
  assign n6253 = ~n3246 ;
  assign n3247 = n3245 & n6253 ;
  assign n6254 = ~n3247 ;
  assign n3254 = x[0] & n6254 ;
  assign n6255 = ~n825 ;
  assign n3260 = n321 & n6255 ;
  assign n6256 = ~n484 ;
  assign n3261 = n6256 & n3260 ;
  assign n6257 = ~n428 ;
  assign n3262 = n6257 & n3261 ;
  assign n6258 = ~n2246 ;
  assign n3263 = n6258 & n3262 ;
  assign n6259 = ~n2336 ;
  assign n3264 = n6259 & n3263 ;
  assign n6260 = ~n2423 ;
  assign n3265 = n6260 & n3264 ;
  assign n6261 = ~n1002 ;
  assign n3266 = n6261 & n3265 ;
  assign n6262 = ~n503 ;
  assign n3267 = n6262 & n3266 ;
  assign n6263 = ~n294 ;
  assign n3268 = n6263 & n3267 ;
  assign n6264 = ~n210 ;
  assign n3269 = n6264 & n3268 ;
  assign n3270 = n5524 & n3269 ;
  assign n6265 = ~n235 ;
  assign n3271 = n6265 & n3270 ;
  assign n3272 = n297 | n824 ;
  assign n3273 = n323 | n3272 ;
  assign n3274 = n198 | n3273 ;
  assign n3275 = n2167 | n3274 ;
  assign n3276 = n412 | n3275 ;
  assign n3277 = n224 | n3276 ;
  assign n3278 = n211 | n3277 ;
  assign n3279 = n367 | n3278 ;
  assign n3280 = n446 | n3279 ;
  assign n3281 = n332 | n3280 ;
  assign n3282 = n110 | n3281 ;
  assign n3283 = n355 | n3282 ;
  assign n3284 = n101 | n3283 ;
  assign n3285 = n339 | n3284 ;
  assign n3286 = n760 | n2370 ;
  assign n3287 = n153 | n3286 ;
  assign n3288 = n784 | n3287 ;
  assign n3289 = n3285 | n3288 ;
  assign n3290 = n208 | n3289 ;
  assign n3291 = n147 | n3290 ;
  assign n3292 = n173 | n3291 ;
  assign n3293 = n218 | n3292 ;
  assign n3294 = n225 | n3293 ;
  assign n3295 = n183 | n3294 ;
  assign n3296 = n445 | n3295 ;
  assign n3297 = n358 | n3296 ;
  assign n3298 = n476 | n3297 ;
  assign n6266 = ~n3298 ;
  assign n3299 = n2556 & n6266 ;
  assign n3300 = n3271 & n3299 ;
  assign n3301 = n131 | n402 ;
  assign n3302 = n346 | n420 ;
  assign n3303 = n1213 | n3302 ;
  assign n3304 = n394 | n3303 ;
  assign n3305 = n434 | n3304 ;
  assign n3306 = n311 | n3305 ;
  assign n3307 = n484 | n3306 ;
  assign n3308 = n501 | n3307 ;
  assign n3309 = n452 | n3308 ;
  assign n3310 = n3301 | n3309 ;
  assign n3311 = n137 | n3310 ;
  assign n3312 = n3300 & n3311 ;
  assign n3313 = n3300 | n3311 ;
  assign n6267 = ~n3312 ;
  assign n3314 = n6267 & n3313 ;
  assign n3317 = n3254 & n3314 ;
  assign n6268 = ~n284 ;
  assign n3324 = n6268 & n3247 ;
  assign n6269 = ~n2556 ;
  assign n3334 = n6269 & n3298 ;
  assign n3335 = n3299 | n3334 ;
  assign n3362 = n3324 & n3335 ;
  assign n3343 = n3271 | n3299 ;
  assign n6270 = ~n3300 ;
  assign n3344 = n6270 & n3343 ;
  assign n6271 = ~x[0] ;
  assign n3354 = n6271 & n3244 ;
  assign n6272 = ~n3344 ;
  assign n3363 = n6272 & n3354 ;
  assign n3364 = n3362 | n3363 ;
  assign n3365 = n3317 | n3364 ;
  assign n3248 = x[0] & n3247 ;
  assign n3345 = n3335 & n6272 ;
  assign n3336 = n2558 & n3335 ;
  assign n3366 = n2676 | n2678 ;
  assign n3367 = n2558 | n3335 ;
  assign n6273 = ~n3336 ;
  assign n3368 = n6273 & n3367 ;
  assign n3370 = n3366 & n3368 ;
  assign n3371 = n3336 | n3370 ;
  assign n6274 = ~n3335 ;
  assign n3352 = n6274 & n3344 ;
  assign n3372 = n3345 | n3352 ;
  assign n6275 = ~n3372 ;
  assign n3374 = n3371 & n6275 ;
  assign n3375 = n3345 | n3374 ;
  assign n3353 = n3314 & n3344 ;
  assign n3376 = n3314 | n3344 ;
  assign n6276 = ~n3353 ;
  assign n3377 = n6276 & n3376 ;
  assign n3378 = n3375 | n3377 ;
  assign n3379 = n3375 & n3377 ;
  assign n6277 = ~n3379 ;
  assign n3380 = n3378 & n6277 ;
  assign n6278 = ~n3380 ;
  assign n3383 = n3248 & n6278 ;
  assign n3384 = n3365 | n3383 ;
  assign n3385 = n5502 & n3384 ;
  assign n6279 = ~n3384 ;
  assign n3386 = n287 & n6279 ;
  assign n3387 = n3385 | n3386 ;
  assign n3388 = n3240 & n3387 ;
  assign n6280 = ~n3234 ;
  assign n3235 = n3086 & n6280 ;
  assign n6281 = ~n3086 ;
  assign n3389 = n6281 & n3234 ;
  assign n3390 = n3235 | n3389 ;
  assign n3346 = n3254 & n6272 ;
  assign n3391 = n2558 & n3324 ;
  assign n3392 = n3335 & n3354 ;
  assign n3393 = n3391 | n3392 ;
  assign n3394 = n3346 | n3393 ;
  assign n3373 = n3371 | n3372 ;
  assign n3395 = n3371 & n3372 ;
  assign n6282 = ~n3395 ;
  assign n3396 = n3373 & n6282 ;
  assign n6283 = ~n3396 ;
  assign n3400 = n3248 & n6283 ;
  assign n3401 = n3394 | n3400 ;
  assign n3402 = n5502 & n3401 ;
  assign n6284 = ~n3401 ;
  assign n3403 = n287 & n6284 ;
  assign n3404 = n3402 | n3403 ;
  assign n3406 = n3390 & n3404 ;
  assign n3326 = n6081 & n3324 ;
  assign n3355 = n2558 & n3354 ;
  assign n3408 = n3326 | n3355 ;
  assign n3409 = n3254 & n3335 ;
  assign n3410 = n3408 | n3409 ;
  assign n6285 = ~n3366 ;
  assign n3369 = n6285 & n3368 ;
  assign n6286 = ~n3368 ;
  assign n3411 = n3366 & n6286 ;
  assign n3412 = n3369 | n3411 ;
  assign n3413 = n3248 & n3412 ;
  assign n3417 = n3410 | n3413 ;
  assign n3418 = n287 | n3417 ;
  assign n3419 = n287 & n3417 ;
  assign n6287 = ~n3419 ;
  assign n3420 = n3418 & n6287 ;
  assign n3428 = n287 & n3248 ;
  assign n3461 = n6145 & n3428 ;
  assign n3429 = n2711 & n3428 ;
  assign n3357 = n2633 & n3354 ;
  assign n6288 = ~n3357 ;
  assign n3466 = n287 & n6288 ;
  assign n3467 = n2630 & n3254 ;
  assign n6289 = ~n3467 ;
  assign n3468 = n3466 & n6289 ;
  assign n6290 = ~n3429 ;
  assign n3469 = n6290 & n3468 ;
  assign n3256 = n6101 & n3254 ;
  assign n3462 = n2633 & n3324 ;
  assign n3463 = n2630 & n3354 ;
  assign n3464 = n3462 | n3463 ;
  assign n3465 = n3256 | n3464 ;
  assign n3470 = n287 & n3465 ;
  assign n6291 = ~n3470 ;
  assign n3471 = n3469 & n6291 ;
  assign n6292 = ~n3461 ;
  assign n3472 = n6292 & n3471 ;
  assign n3473 = x[0] & n2633 ;
  assign n6293 = ~n3473 ;
  assign n3474 = n3472 & n6293 ;
  assign n3475 = n3170 | n3474 ;
  assign n3249 = n6149 & n3248 ;
  assign n3259 = n2616 & n3254 ;
  assign n3329 = n2630 & n3324 ;
  assign n3476 = n3259 | n3329 ;
  assign n3477 = n6101 & n3354 ;
  assign n3478 = n3476 | n3477 ;
  assign n3479 = n3249 | n3478 ;
  assign n3480 = n287 | n3479 ;
  assign n3481 = n287 & n3479 ;
  assign n6294 = ~n3481 ;
  assign n3482 = n3480 & n6294 ;
  assign n3483 = n3475 & n3482 ;
  assign n3484 = n3170 & n3474 ;
  assign n3485 = n3483 | n3484 ;
  assign n3486 = n3171 | n3178 ;
  assign n6295 = ~n3179 ;
  assign n3487 = n6295 & n3486 ;
  assign n3496 = n3485 & n3487 ;
  assign n3325 = n6101 & n3324 ;
  assign n3456 = n2611 & n3254 ;
  assign n3457 = n2616 & n3354 ;
  assign n3458 = n3456 | n3457 ;
  assign n3459 = n3325 | n3458 ;
  assign n3460 = n287 & n3459 ;
  assign n3488 = n3485 | n3487 ;
  assign n3491 = n2760 & n3428 ;
  assign n6296 = ~n3491 ;
  assign n3493 = n3488 & n6296 ;
  assign n3489 = n2760 & n3248 ;
  assign n3490 = n3459 | n3489 ;
  assign n3494 = n287 | n3490 ;
  assign n3495 = n3493 & n3494 ;
  assign n6297 = ~n3460 ;
  assign n3497 = n6297 & n3495 ;
  assign n3498 = n3496 | n3497 ;
  assign n3250 = n2821 & n3248 ;
  assign n3330 = n2616 & n3324 ;
  assign n3358 = n2611 & n3354 ;
  assign n3499 = n3330 | n3358 ;
  assign n3500 = n2605 & n3254 ;
  assign n3501 = n3499 | n3500 ;
  assign n3502 = n3250 | n3501 ;
  assign n3503 = n287 | n3502 ;
  assign n3504 = n287 & n3502 ;
  assign n6298 = ~n3504 ;
  assign n3505 = n3503 & n6298 ;
  assign n3506 = n3498 & n3505 ;
  assign n3455 = n3179 | n3188 ;
  assign n3507 = n3498 | n3505 ;
  assign n6299 = ~n3189 ;
  assign n3508 = n6299 & n3507 ;
  assign n3509 = n3455 & n3508 ;
  assign n3510 = n3506 | n3509 ;
  assign n6300 = ~n3199 ;
  assign n3200 = n3192 & n6300 ;
  assign n6301 = ~n3192 ;
  assign n3511 = n6301 & n3199 ;
  assign n3512 = n3200 | n3511 ;
  assign n3513 = n3510 & n3512 ;
  assign n3255 = n2598 & n3254 ;
  assign n3447 = n2611 & n3324 ;
  assign n3448 = n2605 & n3354 ;
  assign n3449 = n3447 | n3448 ;
  assign n3450 = n3255 | n3449 ;
  assign n3451 = n287 & n3450 ;
  assign n3452 = n2927 & n3248 ;
  assign n3453 = n3450 | n3452 ;
  assign n3454 = n287 | n3453 ;
  assign n3514 = n2927 & n3428 ;
  assign n3515 = n3510 | n3512 ;
  assign n6302 = ~n3514 ;
  assign n3516 = n6302 & n3515 ;
  assign n3517 = n3454 & n3516 ;
  assign n6303 = ~n3451 ;
  assign n3518 = n6303 & n3517 ;
  assign n3519 = n3513 | n3518 ;
  assign n3251 = n6168 & n3248 ;
  assign n3327 = n2605 & n3324 ;
  assign n3359 = n2598 & n3354 ;
  assign n3520 = n3327 | n3359 ;
  assign n3521 = n6091 & n3254 ;
  assign n3522 = n3520 | n3521 ;
  assign n3523 = n3251 | n3522 ;
  assign n3524 = n287 | n3523 ;
  assign n3525 = n287 & n3523 ;
  assign n6304 = ~n3525 ;
  assign n3526 = n3524 & n6304 ;
  assign n3527 = n3519 & n3526 ;
  assign n3446 = n3202 | n3204 ;
  assign n3528 = n3519 | n3526 ;
  assign n6305 = ~n3205 ;
  assign n3529 = n6305 & n3528 ;
  assign n3530 = n3446 & n3529 ;
  assign n3531 = n3527 | n3530 ;
  assign n6306 = ~n3206 ;
  assign n3209 = n6306 & n3208 ;
  assign n6307 = ~n3208 ;
  assign n3532 = n3206 & n6307 ;
  assign n3533 = n3209 | n3532 ;
  assign n3534 = n3531 & n3533 ;
  assign n3258 = n2589 & n3254 ;
  assign n3438 = n2598 & n3324 ;
  assign n3439 = n6091 & n3354 ;
  assign n3440 = n3438 | n3439 ;
  assign n3441 = n3258 | n3440 ;
  assign n3442 = n287 & n3441 ;
  assign n3443 = n6165 & n3248 ;
  assign n3444 = n3441 | n3443 ;
  assign n3445 = n287 | n3444 ;
  assign n3535 = n6165 & n3428 ;
  assign n3536 = n3531 | n3533 ;
  assign n6308 = ~n3535 ;
  assign n3537 = n6308 & n3536 ;
  assign n3538 = n3445 & n3537 ;
  assign n6309 = ~n3442 ;
  assign n3539 = n6309 & n3538 ;
  assign n3540 = n3534 | n3539 ;
  assign n6310 = ~n3212 ;
  assign n3213 = n3211 & n6310 ;
  assign n6311 = ~n3211 ;
  assign n3541 = n6311 & n3212 ;
  assign n3542 = n3213 | n3541 ;
  assign n3543 = n3540 & n3542 ;
  assign n3257 = n2584 & n3254 ;
  assign n3430 = n6091 & n3324 ;
  assign n3431 = n2589 & n3354 ;
  assign n3432 = n3430 | n3431 ;
  assign n3433 = n3257 | n3432 ;
  assign n3434 = n287 & n3433 ;
  assign n3435 = n3051 & n3248 ;
  assign n3436 = n3433 | n3435 ;
  assign n3437 = n287 | n3436 ;
  assign n3544 = n3051 & n3428 ;
  assign n3545 = n3540 | n3542 ;
  assign n6312 = ~n3544 ;
  assign n3546 = n6312 & n3545 ;
  assign n3547 = n3437 & n3546 ;
  assign n6313 = ~n3434 ;
  assign n3548 = n6313 & n3547 ;
  assign n3549 = n3543 | n3548 ;
  assign n6314 = ~n3215 ;
  assign n3218 = n6314 & n3217 ;
  assign n6315 = ~n3217 ;
  assign n3550 = n3215 & n6315 ;
  assign n3551 = n3218 | n3550 ;
  assign n3552 = n3549 & n3551 ;
  assign n3328 = n2589 & n3324 ;
  assign n3356 = n2584 & n3354 ;
  assign n3421 = n3328 | n3356 ;
  assign n3422 = n2564 & n3254 ;
  assign n3423 = n3421 | n3422 ;
  assign n3424 = n287 & n3423 ;
  assign n3425 = n3093 & n3248 ;
  assign n3426 = n3423 | n3425 ;
  assign n3427 = n287 | n3426 ;
  assign n3553 = n3093 & n3428 ;
  assign n3554 = n3549 | n3551 ;
  assign n6316 = ~n3553 ;
  assign n3555 = n6316 & n3554 ;
  assign n3556 = n3427 & n3555 ;
  assign n6317 = ~n3424 ;
  assign n3557 = n6317 & n3556 ;
  assign n3558 = n3552 | n3557 ;
  assign n6318 = ~n3222 ;
  assign n3223 = n3220 & n6318 ;
  assign n6319 = ~n3220 ;
  assign n3559 = n6319 & n3222 ;
  assign n3560 = n3223 | n3559 ;
  assign n3561 = n3558 & n3560 ;
  assign n3252 = n6213 & n3248 ;
  assign n3331 = n2584 & n3324 ;
  assign n3360 = n2564 & n3354 ;
  assign n3562 = n3331 | n3360 ;
  assign n3563 = n6081 & n3254 ;
  assign n3564 = n3562 | n3563 ;
  assign n3565 = n3252 | n3564 ;
  assign n3566 = n287 | n3565 ;
  assign n3567 = n287 & n3565 ;
  assign n6320 = ~n3567 ;
  assign n3568 = n3566 & n6320 ;
  assign n3569 = n3561 | n3568 ;
  assign n3570 = n3558 | n3560 ;
  assign n3571 = n3569 & n3570 ;
  assign n6321 = ~n3227 ;
  assign n3228 = n3225 & n6321 ;
  assign n6322 = ~n3225 ;
  assign n3572 = n6322 & n3227 ;
  assign n3573 = n3228 | n3572 ;
  assign n3574 = n3571 | n3573 ;
  assign n3253 = n6124 & n3248 ;
  assign n3332 = n2564 & n3324 ;
  assign n3361 = n6081 & n3354 ;
  assign n3575 = n3332 | n3361 ;
  assign n3576 = n2558 & n3254 ;
  assign n3577 = n3575 | n3576 ;
  assign n3578 = n3253 | n3577 ;
  assign n3579 = n287 | n3578 ;
  assign n3580 = n287 & n3578 ;
  assign n6323 = ~n3580 ;
  assign n3581 = n3579 & n6323 ;
  assign n3582 = n3574 & n3581 ;
  assign n3583 = n3571 & n3573 ;
  assign n3584 = n3582 | n3583 ;
  assign n3585 = n3420 & n3584 ;
  assign n3407 = n3230 | n3232 ;
  assign n3586 = n3420 | n3584 ;
  assign n6324 = ~n3233 ;
  assign n3587 = n6324 & n3586 ;
  assign n3588 = n3407 & n3587 ;
  assign n3589 = n3585 | n3588 ;
  assign n6325 = ~n3390 ;
  assign n3405 = n6325 & n3404 ;
  assign n6326 = ~n3404 ;
  assign n3590 = n3390 & n6326 ;
  assign n3591 = n3405 | n3590 ;
  assign n3592 = n3589 & n3591 ;
  assign n3593 = n3406 | n3592 ;
  assign n6327 = ~n3387 ;
  assign n3594 = n3240 & n6327 ;
  assign n6328 = ~n3240 ;
  assign n3595 = n6328 & n3387 ;
  assign n3596 = n3594 | n3595 ;
  assign n3597 = n3593 & n3596 ;
  assign n3598 = n3388 | n3597 ;
  assign n3599 = n3070 & n3237 ;
  assign n3600 = n3069 | n3599 ;
  assign n3414 = n2581 & n3412 ;
  assign n2571 = n2562 & n6081 ;
  assign n2577 = n2558 & n2574 ;
  assign n3601 = n2571 | n2577 ;
  assign n3602 = n292 & n3335 ;
  assign n3603 = n3601 | n3602 ;
  assign n3604 = n3414 | n3603 ;
  assign n6329 = ~n3604 ;
  assign n3605 = n274 & n6329 ;
  assign n3606 = n5721 & n3604 ;
  assign n3607 = n3605 | n3606 ;
  assign n3062 = n3049 & n3060 ;
  assign n3608 = n3017 & n3064 ;
  assign n3609 = n3062 | n3608 ;
  assign n3610 = n3025 & n3041 ;
  assign n3611 = n3048 | n3610 ;
  assign n2911 = n2727 & n6168 ;
  assign n2737 = n2605 & n2733 ;
  assign n2745 = n2598 & n2742 ;
  assign n3612 = n2737 | n2745 ;
  assign n3613 = n6091 & n2748 ;
  assign n3614 = n3612 | n3613 ;
  assign n3615 = n2911 | n3614 ;
  assign n6330 = ~n3615 ;
  assign n3616 = n672 & n6330 ;
  assign n3617 = n5514 & n3615 ;
  assign n3618 = n3616 | n3617 ;
  assign n3619 = n523 & n2630 ;
  assign n3492 = n2713 & n2760 ;
  assign n2694 = n2616 & n2693 ;
  assign n2702 = n2611 & n2699 ;
  assign n3620 = n2694 | n2702 ;
  assign n3621 = n6101 & n2831 ;
  assign n3622 = n3620 | n3621 ;
  assign n3623 = n3492 | n3622 ;
  assign n3625 = n523 & n3623 ;
  assign n6331 = ~n3625 ;
  assign n3626 = n3619 & n6331 ;
  assign n6332 = ~n3623 ;
  assign n3624 = n523 & n6332 ;
  assign n3627 = n5542 & n3623 ;
  assign n3628 = n3624 | n3627 ;
  assign n3629 = n3619 | n3628 ;
  assign n6333 = ~n3626 ;
  assign n3630 = n6333 & n3629 ;
  assign n6334 = ~n3630 ;
  assign n3631 = n3039 & n6334 ;
  assign n3632 = n6198 & n3630 ;
  assign n3633 = n3631 | n3632 ;
  assign n6335 = ~n3633 ;
  assign n3634 = n3618 & n6335 ;
  assign n6336 = ~n3618 ;
  assign n3635 = n6336 & n3633 ;
  assign n3636 = n3634 | n3635 ;
  assign n3637 = n3611 | n3636 ;
  assign n3638 = n3611 & n3636 ;
  assign n6337 = ~n3638 ;
  assign n3639 = n3637 & n6337 ;
  assign n2866 = n2564 & n2860 ;
  assign n3640 = n2589 & n2870 ;
  assign n3641 = n2584 & n2879 ;
  assign n3642 = n3640 | n3641 ;
  assign n3643 = n2866 | n3642 ;
  assign n3644 = n2891 & n3093 ;
  assign n3645 = n3643 | n3644 ;
  assign n3646 = n1052 & n3645 ;
  assign n3647 = n1052 | n3645 ;
  assign n6338 = ~n3646 ;
  assign n3648 = n6338 & n3647 ;
  assign n3649 = n3639 & n3648 ;
  assign n3650 = n3639 | n3648 ;
  assign n6339 = ~n3649 ;
  assign n3651 = n6339 & n3650 ;
  assign n6340 = ~n3609 ;
  assign n3652 = n6340 & n3651 ;
  assign n6341 = ~n3651 ;
  assign n3653 = n3609 & n6341 ;
  assign n3654 = n3652 | n3653 ;
  assign n3655 = n3607 & n3654 ;
  assign n3656 = n3607 | n3654 ;
  assign n6342 = ~n3655 ;
  assign n3657 = n6342 & n3656 ;
  assign n6343 = ~n3600 ;
  assign n3658 = n6343 & n3657 ;
  assign n6344 = ~n3657 ;
  assign n3659 = n3600 & n6344 ;
  assign n3660 = n3658 | n3659 ;
  assign n3661 = n345 | n501 ;
  assign n3662 = n145 | n3661 ;
  assign n3663 = n513 | n3662 ;
  assign n3664 = n484 | n3663 ;
  assign n3665 = n411 | n3664 ;
  assign n3666 = n401 | n3665 ;
  assign n3667 = n186 | n3666 ;
  assign n3668 = n217 | n3667 ;
  assign n3669 = n222 | n3668 ;
  assign n6345 = ~n3311 ;
  assign n3670 = n3300 & n6345 ;
  assign n6346 = ~n3669 ;
  assign n3671 = n6346 & n3670 ;
  assign n6347 = ~n3670 ;
  assign n3672 = n3669 & n6347 ;
  assign n3673 = n3671 | n3672 ;
  assign n3674 = n3254 & n3673 ;
  assign n3685 = n3324 & n6272 ;
  assign n3686 = n3314 & n3354 ;
  assign n3687 = n3685 | n3686 ;
  assign n3688 = n3674 | n3687 ;
  assign n3689 = n3314 & n6272 ;
  assign n6348 = ~n3377 ;
  assign n3690 = n3375 & n6348 ;
  assign n3691 = n3689 | n3690 ;
  assign n6349 = ~n3673 ;
  assign n3684 = n3314 & n6349 ;
  assign n6350 = ~n3314 ;
  assign n3692 = n6350 & n3673 ;
  assign n3693 = n3684 | n3692 ;
  assign n6351 = ~n3691 ;
  assign n3694 = n6351 & n3693 ;
  assign n6352 = ~n3693 ;
  assign n3695 = n3691 & n6352 ;
  assign n3696 = n3694 | n3695 ;
  assign n3699 = n3248 & n3696 ;
  assign n3700 = n3688 | n3699 ;
  assign n3701 = n5502 & n3700 ;
  assign n6353 = ~n3700 ;
  assign n3702 = n287 & n6353 ;
  assign n3703 = n3701 | n3702 ;
  assign n3704 = n3660 & n3703 ;
  assign n3705 = n3660 | n3703 ;
  assign n6354 = ~n3704 ;
  assign n3706 = n6354 & n3705 ;
  assign n6355 = ~n3598 ;
  assign n3707 = n6355 & n3706 ;
  assign n6356 = ~n3706 ;
  assign n3708 = n3598 & n6356 ;
  assign n3709 = n3707 | n3708 ;
  assign n3711 = n269 & n3709 ;
  assign n3710 = n269 | n3709 ;
  assign n6357 = ~n3711 ;
  assign n3781 = n3710 & n6357 ;
  assign n3712 = n110 | n505 ;
  assign n3713 = n752 | n3712 ;
  assign n3714 = n293 | n3713 ;
  assign n3715 = n151 | n3714 ;
  assign n3716 = n822 | n3715 ;
  assign n3717 = n136 | n3716 ;
  assign n3718 = n147 | n3717 ;
  assign n3719 = n183 | n3718 ;
  assign n3720 = n310 | n3719 ;
  assign n3721 = n130 | n3720 ;
  assign n3722 = n356 | n3721 ;
  assign n3723 = n139 | n3722 ;
  assign n3724 = n101 | n3723 ;
  assign n3725 = n369 | n504 ;
  assign n3726 = n1182 | n3725 ;
  assign n3727 = n215 | n3726 ;
  assign n3728 = n253 | n3727 ;
  assign n3729 = n494 | n3728 ;
  assign n3730 = n552 | n3729 ;
  assign n3731 = n444 | n3730 ;
  assign n3732 = n470 | n3731 ;
  assign n3733 = n213 | n3732 ;
  assign n3734 = n805 | n3733 ;
  assign n3735 = n414 | n3734 ;
  assign n3736 = n295 | n3735 ;
  assign n3737 = n2459 | n3736 ;
  assign n3738 = n3724 | n3737 ;
  assign n3739 = n1006 | n3738 ;
  assign n3740 = n134 | n3739 ;
  assign n3741 = n252 | n3740 ;
  assign n3742 = n324 | n3741 ;
  assign n3743 = n445 | n3742 ;
  assign n3744 = n143 | n3743 ;
  assign n3745 = n294 | n3744 ;
  assign n3746 = n332 | n3745 ;
  assign n3747 = n469 | n3746 ;
  assign n3748 = n339 | n3747 ;
  assign n3750 = n3593 | n3595 ;
  assign n3751 = n3594 | n3750 ;
  assign n6358 = ~n3597 ;
  assign n3752 = n6358 & n3751 ;
  assign n3753 = n394 | n2280 ;
  assign n3754 = n2306 | n3753 ;
  assign n3755 = n141 | n3754 ;
  assign n3756 = n502 | n3755 ;
  assign n3757 = n353 | n3756 ;
  assign n3758 = n476 | n3757 ;
  assign n3759 = n338 | n829 ;
  assign n3760 = n134 | n3759 ;
  assign n3761 = n152 | n3760 ;
  assign n3762 = n459 | n2427 ;
  assign n3763 = n2438 | n3762 ;
  assign n3764 = n341 | n3763 ;
  assign n3765 = n3761 | n3764 ;
  assign n3766 = n3758 | n3765 ;
  assign n3767 = n2368 | n3766 ;
  assign n3768 = n412 | n3767 ;
  assign n3769 = n147 | n3768 ;
  assign n3770 = n314 | n3769 ;
  assign n3771 = n217 | n3770 ;
  assign n3772 = n171 | n3771 ;
  assign n3773 = n216 | n3772 ;
  assign n3774 = n299 | n3773 ;
  assign n6359 = ~n3591 ;
  assign n3749 = n3589 & n6359 ;
  assign n6360 = ~n3589 ;
  assign n3775 = n6360 & n3591 ;
  assign n3776 = n3749 | n3775 ;
  assign n3777 = n3774 & n3776 ;
  assign n3778 = n3752 | n3777 ;
  assign n3779 = n3748 & n3778 ;
  assign n3780 = n3752 & n3777 ;
  assign n3782 = n3779 | n3780 ;
  assign n3783 = n3781 & n3782 ;
  assign n3784 = n3711 | n3783 ;
  assign n3333 = n3314 & n3324 ;
  assign n3675 = n3354 & n3673 ;
  assign n3814 = n3333 | n3675 ;
  assign n3785 = n237 | n589 ;
  assign n3786 = n347 | n3785 ;
  assign n3787 = n120 | n3786 ;
  assign n3788 = n310 | n3787 ;
  assign n3789 = n205 | n3788 ;
  assign n3790 = n444 | n3789 ;
  assign n3791 = n468 | n3790 ;
  assign n3792 = n350 | n467 ;
  assign n3793 = n331 | n3792 ;
  assign n6361 = ~n3793 ;
  assign n3794 = n1210 & n6361 ;
  assign n6362 = ~n3791 ;
  assign n3795 = n6362 & n3794 ;
  assign n3796 = n6260 & n3795 ;
  assign n6363 = ~n220 ;
  assign n3797 = n6363 & n3796 ;
  assign n6364 = ~n314 ;
  assign n3798 = n6364 & n3797 ;
  assign n6365 = ~n174 ;
  assign n3799 = n6365 & n3798 ;
  assign n6366 = ~n216 ;
  assign n3800 = n6366 & n3799 ;
  assign n6367 = ~n553 ;
  assign n3801 = n6367 & n3800 ;
  assign n3802 = n5741 & n3801 ;
  assign n6368 = ~n129 ;
  assign n3803 = n6368 & n3802 ;
  assign n6369 = ~n221 ;
  assign n3804 = n6369 & n3803 ;
  assign n6370 = ~n3804 ;
  assign n3805 = n3671 & n6370 ;
  assign n6371 = ~n3671 ;
  assign n3806 = n6371 & n3804 ;
  assign n3807 = n3805 | n3806 ;
  assign n6372 = ~n3807 ;
  assign n3815 = n3254 & n6372 ;
  assign n3816 = n3814 | n3815 ;
  assign n3817 = n3314 & n3673 ;
  assign n3818 = n3691 & n3693 ;
  assign n3819 = n3817 | n3818 ;
  assign n3809 = n3673 & n6372 ;
  assign n3820 = n6349 & n3807 ;
  assign n3821 = n3809 | n3820 ;
  assign n6373 = ~n3819 ;
  assign n3822 = n6373 & n3821 ;
  assign n6374 = ~n3821 ;
  assign n3823 = n3819 & n6374 ;
  assign n3824 = n3822 | n3823 ;
  assign n6375 = ~n3824 ;
  assign n3825 = n3248 & n6375 ;
  assign n3829 = n3816 | n3825 ;
  assign n3830 = n287 | n3829 ;
  assign n3831 = n287 & n3829 ;
  assign n6376 = ~n3831 ;
  assign n3832 = n3830 & n6376 ;
  assign n3833 = n3600 & n3657 ;
  assign n3834 = n3655 | n3833 ;
  assign n3079 = n2891 & n6213 ;
  assign n2875 = n2584 & n2870 ;
  assign n2883 = n2564 & n2879 ;
  assign n3835 = n2875 | n2883 ;
  assign n3836 = n6081 & n2860 ;
  assign n3837 = n3835 | n3836 ;
  assign n3838 = n3079 | n3837 ;
  assign n6377 = ~n3838 ;
  assign n3839 = n1052 & n6377 ;
  assign n3840 = n5595 & n3838 ;
  assign n3841 = n3839 | n3840 ;
  assign n3842 = n3618 & n3633 ;
  assign n3843 = n3638 | n3842 ;
  assign n3844 = n3039 & n3630 ;
  assign n3845 = n3626 | n3844 ;
  assign n2824 = n2713 & n2821 ;
  assign n2695 = n2611 & n2693 ;
  assign n2833 = n2616 & n2831 ;
  assign n3846 = n2695 | n2833 ;
  assign n3847 = n2605 & n2699 ;
  assign n3848 = n3846 | n3847 ;
  assign n3849 = n2824 | n3848 ;
  assign n3851 = n523 & n2624 ;
  assign n6378 = ~n3849 ;
  assign n3852 = n6378 & n3851 ;
  assign n6379 = ~n3851 ;
  assign n3853 = n3849 & n6379 ;
  assign n3854 = n3852 | n3853 ;
  assign n6380 = ~n3845 ;
  assign n3855 = n6380 & n3854 ;
  assign n6381 = ~n3854 ;
  assign n3856 = n3845 & n6381 ;
  assign n3857 = n3855 | n3856 ;
  assign n2749 = n2589 & n2748 ;
  assign n3858 = n2598 & n2733 ;
  assign n3859 = n6091 & n2742 ;
  assign n3860 = n3858 | n3859 ;
  assign n3861 = n2749 | n3860 ;
  assign n3862 = n2727 & n6165 ;
  assign n3863 = n3861 | n3862 ;
  assign n3864 = n672 & n3863 ;
  assign n3865 = n672 | n3863 ;
  assign n6382 = ~n3864 ;
  assign n3866 = n6382 & n3865 ;
  assign n6383 = ~n3857 ;
  assign n3867 = n6383 & n3866 ;
  assign n6384 = ~n3866 ;
  assign n3868 = n3857 & n6384 ;
  assign n3869 = n3867 | n3868 ;
  assign n6385 = ~n3869 ;
  assign n3870 = n3843 & n6385 ;
  assign n6386 = ~n3843 ;
  assign n3871 = n6386 & n3869 ;
  assign n3872 = n3870 | n3871 ;
  assign n3873 = n3841 | n3872 ;
  assign n3874 = n3841 & n3872 ;
  assign n6387 = ~n3874 ;
  assign n3875 = n3873 & n6387 ;
  assign n3876 = n3609 & n3651 ;
  assign n3877 = n3649 | n3876 ;
  assign n3878 = n3875 | n3877 ;
  assign n3879 = n3875 & n3877 ;
  assign n6388 = ~n3879 ;
  assign n3880 = n3878 & n6388 ;
  assign n3347 = n292 & n6272 ;
  assign n3881 = n2558 & n2562 ;
  assign n3882 = n2574 & n3335 ;
  assign n3883 = n3881 | n3882 ;
  assign n3884 = n3347 | n3883 ;
  assign n3885 = n2581 & n6283 ;
  assign n3886 = n3884 | n3885 ;
  assign n3887 = n274 & n3886 ;
  assign n3888 = n274 | n3886 ;
  assign n6389 = ~n3887 ;
  assign n3889 = n6389 & n3888 ;
  assign n6390 = ~n3880 ;
  assign n3890 = n6390 & n3889 ;
  assign n6391 = ~n3889 ;
  assign n3891 = n3880 & n6391 ;
  assign n3892 = n3890 | n3891 ;
  assign n6392 = ~n3892 ;
  assign n3893 = n3834 & n6392 ;
  assign n6393 = ~n3834 ;
  assign n3894 = n6393 & n3892 ;
  assign n3895 = n3893 | n3894 ;
  assign n6394 = ~n3895 ;
  assign n3896 = n3832 & n6394 ;
  assign n6395 = ~n3832 ;
  assign n3897 = n6395 & n3895 ;
  assign n3898 = n3896 | n3897 ;
  assign n3899 = n3598 & n3706 ;
  assign n3900 = n3704 | n3899 ;
  assign n3901 = n3898 | n3900 ;
  assign n3902 = n3898 & n3900 ;
  assign n6396 = ~n3902 ;
  assign n3903 = n3901 & n6396 ;
  assign n3904 = n237 | n1140 ;
  assign n3905 = n822 | n3904 ;
  assign n3906 = n1516 | n3905 ;
  assign n3907 = n2314 | n3906 ;
  assign n3908 = n642 | n3907 ;
  assign n3909 = n622 | n3908 ;
  assign n3910 = n208 | n3909 ;
  assign n3911 = n253 | n3910 ;
  assign n3912 = n145 | n3911 ;
  assign n3913 = n342 | n3912 ;
  assign n6397 = ~n3913 ;
  assign n3914 = n3903 & n6397 ;
  assign n6398 = ~n3903 ;
  assign n3915 = n6398 & n3913 ;
  assign n3916 = n3914 | n3915 ;
  assign n3917 = n3784 | n3916 ;
  assign n3918 = n3784 & n3916 ;
  assign n6399 = ~n3918 ;
  assign n3919 = n3917 & n6399 ;
  assign n3920 = n3781 | n3782 ;
  assign n6400 = ~n3783 ;
  assign n3921 = n6400 & n3920 ;
  assign n3922 = n3919 | n3921 ;
  assign n3923 = n3919 & n3921 ;
  assign n6401 = ~n3923 ;
  assign n25 = n3922 & n6401 ;
  assign n3925 = n3903 & n3913 ;
  assign n3926 = n3918 | n3925 ;
  assign n3676 = n3324 & n3673 ;
  assign n3810 = n3354 & n6372 ;
  assign n3957 = n3676 | n3810 ;
  assign n3927 = n3671 & n3804 ;
  assign n3928 = n234 | n2438 ;
  assign n3929 = n456 | n3928 ;
  assign n3930 = n769 | n3929 ;
  assign n3931 = n166 | n3930 ;
  assign n3932 = n114 | n3931 ;
  assign n3933 = n163 | n3932 ;
  assign n3934 = n165 | n3933 ;
  assign n3935 = n313 | n554 ;
  assign n3936 = n831 | n3935 ;
  assign n6402 = ~n3936 ;
  assign n3937 = n1533 & n6402 ;
  assign n6403 = ~n3934 ;
  assign n3938 = n6403 & n3937 ;
  assign n3939 = n6029 & n3938 ;
  assign n3940 = n6261 & n3939 ;
  assign n6404 = ~n494 ;
  assign n3941 = n6404 & n3940 ;
  assign n6405 = ~n469 ;
  assign n3942 = n6405 & n3941 ;
  assign n6406 = ~n364 ;
  assign n3943 = n6406 & n3942 ;
  assign n6407 = ~n323 ;
  assign n3944 = n6407 & n3943 ;
  assign n3945 = n3927 & n3944 ;
  assign n3946 = n3927 | n3944 ;
  assign n6408 = ~n3945 ;
  assign n3947 = n6408 & n3946 ;
  assign n6409 = ~n3947 ;
  assign n3958 = n3254 & n6409 ;
  assign n3959 = n3957 | n3958 ;
  assign n3960 = n3809 | n3823 ;
  assign n3950 = n3807 & n6409 ;
  assign n3961 = n6372 & n3947 ;
  assign n3962 = n3950 | n3961 ;
  assign n3963 = n3960 & n3962 ;
  assign n3964 = n3960 | n3962 ;
  assign n6410 = ~n3963 ;
  assign n3965 = n6410 & n3964 ;
  assign n3966 = n3248 & n3965 ;
  assign n3969 = n3959 | n3966 ;
  assign n3970 = n287 | n3969 ;
  assign n3971 = n287 & n3969 ;
  assign n6411 = ~n3971 ;
  assign n3972 = n3970 & n6411 ;
  assign n3973 = n3880 & n3889 ;
  assign n3974 = n3834 & n3892 ;
  assign n3975 = n3973 | n3974 ;
  assign n2892 = n6124 & n2891 ;
  assign n2876 = n2564 & n2870 ;
  assign n2884 = n6081 & n2879 ;
  assign n3976 = n2876 | n2884 ;
  assign n3977 = n2558 & n2860 ;
  assign n3978 = n3976 | n3977 ;
  assign n3979 = n2892 | n3978 ;
  assign n6412 = ~n3979 ;
  assign n3980 = n1052 & n6412 ;
  assign n3981 = n5595 & n3979 ;
  assign n3982 = n3980 | n3981 ;
  assign n3983 = n3857 & n3866 ;
  assign n3984 = n3843 & n3869 ;
  assign n3985 = n3983 | n3984 ;
  assign n2626 = n523 & n6101 ;
  assign n3850 = n2626 & n6378 ;
  assign n3986 = n3845 & n3854 ;
  assign n3987 = n3850 | n3986 ;
  assign n2703 = n2598 & n2699 ;
  assign n3988 = n2605 & n2693 ;
  assign n3989 = n2611 & n2831 ;
  assign n3990 = n3988 | n3989 ;
  assign n3991 = n2703 | n3990 ;
  assign n3992 = n2713 & n2927 ;
  assign n3993 = n3991 | n3992 ;
  assign n3994 = n523 & n6107 ;
  assign n3995 = n3993 & n3994 ;
  assign n3996 = n3993 | n3994 ;
  assign n6413 = ~n3995 ;
  assign n3997 = n6413 & n3996 ;
  assign n6414 = ~n3987 ;
  assign n3998 = n6414 & n3997 ;
  assign n6415 = ~n3997 ;
  assign n3999 = n3987 & n6415 ;
  assign n4000 = n3998 | n3999 ;
  assign n2753 = n2584 & n2748 ;
  assign n4001 = n6091 & n2733 ;
  assign n4002 = n2589 & n2742 ;
  assign n4003 = n4001 | n4002 ;
  assign n4004 = n2753 | n4003 ;
  assign n4005 = n2727 & n3051 ;
  assign n4006 = n4004 | n4005 ;
  assign n4007 = n672 & n4006 ;
  assign n4008 = n672 | n4006 ;
  assign n6416 = ~n4007 ;
  assign n4009 = n6416 & n4008 ;
  assign n6417 = ~n4000 ;
  assign n4010 = n6417 & n4009 ;
  assign n6418 = ~n4009 ;
  assign n4011 = n4000 & n6418 ;
  assign n4012 = n4010 | n4011 ;
  assign n6419 = ~n4012 ;
  assign n4013 = n3985 & n6419 ;
  assign n6420 = ~n3985 ;
  assign n4014 = n6420 & n4012 ;
  assign n4015 = n4013 | n4014 ;
  assign n4016 = n3982 | n4015 ;
  assign n4017 = n3982 & n4015 ;
  assign n6421 = ~n4017 ;
  assign n4018 = n4016 & n6421 ;
  assign n4019 = n3874 | n3879 ;
  assign n4020 = n4018 | n4019 ;
  assign n4021 = n4018 & n4019 ;
  assign n6422 = ~n4021 ;
  assign n4022 = n4020 & n6422 ;
  assign n3319 = n292 & n3314 ;
  assign n4023 = n2562 & n3335 ;
  assign n4024 = n2574 & n6272 ;
  assign n4025 = n4023 | n4024 ;
  assign n4026 = n3319 | n4025 ;
  assign n4027 = n2581 & n6278 ;
  assign n4028 = n4026 | n4027 ;
  assign n4029 = n274 & n4028 ;
  assign n4030 = n274 | n4028 ;
  assign n6423 = ~n4029 ;
  assign n4031 = n6423 & n4030 ;
  assign n6424 = ~n4022 ;
  assign n4032 = n6424 & n4031 ;
  assign n6425 = ~n4031 ;
  assign n4033 = n4022 & n6425 ;
  assign n4034 = n4032 | n4033 ;
  assign n6426 = ~n4034 ;
  assign n4035 = n3975 & n6426 ;
  assign n6427 = ~n3975 ;
  assign n4036 = n6427 & n4034 ;
  assign n4037 = n4035 | n4036 ;
  assign n4038 = n3972 | n4037 ;
  assign n4039 = n3972 & n4037 ;
  assign n6428 = ~n4039 ;
  assign n4040 = n4038 & n6428 ;
  assign n4041 = n3832 & n3895 ;
  assign n4042 = n3832 | n3895 ;
  assign n6429 = ~n4041 ;
  assign n4043 = n6429 & n4042 ;
  assign n4044 = n3598 & n3705 ;
  assign n4045 = n3704 | n4044 ;
  assign n4046 = n4043 & n4045 ;
  assign n4047 = n4041 | n4046 ;
  assign n6430 = ~n4047 ;
  assign n4048 = n4040 & n6430 ;
  assign n6431 = ~n4040 ;
  assign n4049 = n6431 & n4047 ;
  assign n4050 = n4048 | n4049 ;
  assign n4051 = n137 | n402 ;
  assign n4052 = n358 | n4051 ;
  assign n4053 = n256 | n4052 ;
  assign n4054 = n636 | n2343 ;
  assign n4055 = n2278 | n4054 ;
  assign n4056 = n247 | n4055 ;
  assign n4057 = n769 | n4056 ;
  assign n4058 = n4053 | n4057 ;
  assign n4059 = n208 | n4058 ;
  assign n4060 = n3273 | n4059 ;
  assign n4061 = n172 | n4060 ;
  assign n4062 = n152 | n4061 ;
  assign n4063 = n324 | n4062 ;
  assign n4064 = n189 | n4063 ;
  assign n4065 = n114 | n4064 ;
  assign n4066 = n444 | n4065 ;
  assign n4067 = n4050 | n4066 ;
  assign n4068 = n4050 & n4066 ;
  assign n6432 = ~n4068 ;
  assign n4069 = n4067 & n6432 ;
  assign n4070 = n3926 & n4069 ;
  assign n4071 = n3926 | n4069 ;
  assign n6433 = ~n4070 ;
  assign n4072 = n6433 & n4071 ;
  assign n4073 = n3923 & n4072 ;
  assign n4074 = n3923 | n4072 ;
  assign n6434 = ~n4073 ;
  assign n4075 = n6434 & n4074 ;
  assign n5176 = x[22] & x[23] ;
  assign n4076 = x[22] | x[23] ;
  assign n6435 = ~n5176 ;
  assign n4077 = n6435 & n4076 ;
  assign n4078 = n25 & n4077 ;
  assign n4079 = n4075 & n4078 ;
  assign n4080 = n4075 | n4078 ;
  assign n6436 = ~n4079 ;
  assign n26 = n6436 & n4080 ;
  assign n4082 = n4068 | n4070 ;
  assign n4083 = n343 | n405 ;
  assign n4084 = n126 | n4083 ;
  assign n4085 = n226 | n4084 ;
  assign n4086 = n139 | n4085 ;
  assign n4087 = n129 | n4086 ;
  assign n4088 = n413 | n607 ;
  assign n4089 = n821 | n4088 ;
  assign n4090 = n4087 | n4089 ;
  assign n4091 = n3758 | n4090 ;
  assign n4092 = n310 | n4091 ;
  assign n4093 = n457 | n4092 ;
  assign n4094 = n503 | n4093 ;
  assign n4095 = n295 | n4094 ;
  assign n4096 = n143 | n4095 ;
  assign n4097 = n505 | n4096 ;
  assign n4098 = n323 | n4097 ;
  assign n6437 = ~n4037 ;
  assign n4099 = n3972 & n6437 ;
  assign n6438 = ~n3972 ;
  assign n4100 = n6438 & n4037 ;
  assign n4101 = n4099 | n4100 ;
  assign n4102 = n4047 & n4101 ;
  assign n4103 = n4039 | n4102 ;
  assign n4104 = n3324 & n6372 ;
  assign n4105 = n3354 & n6409 ;
  assign n4106 = n4104 | n4105 ;
  assign n4108 = n3947 & n6410 ;
  assign n4107 = n3807 & n6410 ;
  assign n4109 = n3947 | n4107 ;
  assign n6439 = ~n4108 ;
  assign n4115 = n6439 & n4109 ;
  assign n4116 = n3248 & n4115 ;
  assign n4120 = n4106 | n4116 ;
  assign n4121 = n287 | n4120 ;
  assign n4123 = n287 & n4120 ;
  assign n6440 = ~n4123 ;
  assign n4124 = n4121 & n6440 ;
  assign n4125 = n4022 & n4031 ;
  assign n4126 = n3975 & n4034 ;
  assign n4127 = n4125 | n4126 ;
  assign n3415 = n2891 & n3412 ;
  assign n2877 = n6081 & n2870 ;
  assign n2881 = n2558 & n2879 ;
  assign n4128 = n2877 | n2881 ;
  assign n4129 = n2860 & n3335 ;
  assign n4130 = n4128 | n4129 ;
  assign n4131 = n3415 | n4130 ;
  assign n6441 = ~n4131 ;
  assign n4132 = n1052 & n6441 ;
  assign n4133 = n5595 & n4131 ;
  assign n4134 = n4132 | n4133 ;
  assign n4135 = n4000 & n4009 ;
  assign n4136 = n3985 & n4012 ;
  assign n4137 = n4135 | n4136 ;
  assign n4138 = n3987 & n3997 ;
  assign n6442 = ~n3993 ;
  assign n4139 = n523 & n6442 ;
  assign n4140 = n2616 & n4139 ;
  assign n4141 = n4138 | n4140 ;
  assign n2909 = n2713 & n6168 ;
  assign n2704 = n6091 & n2699 ;
  assign n4142 = n2598 & n2693 ;
  assign n4143 = n2605 & n2831 ;
  assign n4144 = n4142 | n4143 ;
  assign n4145 = n2704 | n4144 ;
  assign n4146 = n2909 | n4145 ;
  assign n4147 = n523 & n6110 ;
  assign n4148 = n4146 & n4147 ;
  assign n4149 = n4146 | n4147 ;
  assign n6443 = ~n4148 ;
  assign n4150 = n6443 & n4149 ;
  assign n6444 = ~n4141 ;
  assign n4151 = n6444 & n4150 ;
  assign n6445 = ~n4150 ;
  assign n4152 = n4141 & n6445 ;
  assign n4153 = n4151 | n4152 ;
  assign n2754 = n2564 & n2748 ;
  assign n4154 = n2589 & n2733 ;
  assign n4155 = n2584 & n2742 ;
  assign n4156 = n4154 | n4155 ;
  assign n4157 = n2754 | n4156 ;
  assign n4158 = n2727 & n3093 ;
  assign n4159 = n4157 | n4158 ;
  assign n4160 = n672 & n4159 ;
  assign n4161 = n672 | n4159 ;
  assign n6446 = ~n4160 ;
  assign n4162 = n6446 & n4161 ;
  assign n6447 = ~n4153 ;
  assign n4163 = n6447 & n4162 ;
  assign n6448 = ~n4162 ;
  assign n4164 = n4153 & n6448 ;
  assign n4165 = n4163 | n4164 ;
  assign n6449 = ~n4165 ;
  assign n4166 = n4137 & n6449 ;
  assign n6450 = ~n4137 ;
  assign n4167 = n6450 & n4165 ;
  assign n4168 = n4166 | n4167 ;
  assign n4169 = n4134 | n4168 ;
  assign n4170 = n4134 & n4168 ;
  assign n6451 = ~n4170 ;
  assign n4171 = n4169 & n6451 ;
  assign n4172 = n4017 | n4021 ;
  assign n4173 = n4171 | n4172 ;
  assign n4174 = n4171 & n4172 ;
  assign n6452 = ~n4174 ;
  assign n4175 = n4173 & n6452 ;
  assign n3677 = n292 & n3673 ;
  assign n4176 = n2574 & n3314 ;
  assign n4177 = n2562 & n6272 ;
  assign n4178 = n4176 | n4177 ;
  assign n4179 = n3677 | n4178 ;
  assign n4180 = n2581 & n3696 ;
  assign n4181 = n4179 | n4180 ;
  assign n4182 = n274 & n4181 ;
  assign n4183 = n274 | n4181 ;
  assign n6453 = ~n4182 ;
  assign n4184 = n6453 & n4183 ;
  assign n6454 = ~n4184 ;
  assign n4185 = n4175 & n6454 ;
  assign n6455 = ~n4175 ;
  assign n4186 = n6455 & n4184 ;
  assign n4187 = n4185 | n4186 ;
  assign n6456 = ~n4187 ;
  assign n4188 = n4127 & n6456 ;
  assign n6457 = ~n4127 ;
  assign n4189 = n6457 & n4187 ;
  assign n4190 = n4188 | n4189 ;
  assign n6458 = ~n4190 ;
  assign n4191 = n4124 & n6458 ;
  assign n6459 = ~n4124 ;
  assign n4192 = n6459 & n4190 ;
  assign n4193 = n4191 | n4192 ;
  assign n6460 = ~n4193 ;
  assign n4194 = n4103 & n6460 ;
  assign n6461 = ~n4103 ;
  assign n4195 = n6461 & n4193 ;
  assign n4196 = n4194 | n4195 ;
  assign n4198 = n4098 & n4196 ;
  assign n4197 = n4098 | n4196 ;
  assign n4199 = n4082 & n4197 ;
  assign n6462 = ~n4198 ;
  assign n4200 = n6462 & n4199 ;
  assign n6463 = ~n4200 ;
  assign n4201 = n4082 & n6463 ;
  assign n4202 = n4198 | n4199 ;
  assign n6464 = ~n4202 ;
  assign n4203 = n4197 & n6464 ;
  assign n4204 = n4201 | n4203 ;
  assign n4205 = n4073 | n4204 ;
  assign n4206 = n4073 & n4204 ;
  assign n6465 = ~n4206 ;
  assign n4207 = n4205 & n6465 ;
  assign n4208 = n25 | n4075 ;
  assign n4209 = n4077 & n4208 ;
  assign n4210 = n4207 & n4209 ;
  assign n4211 = n4207 | n4209 ;
  assign n6466 = ~n4210 ;
  assign n27 = n6466 & n4211 ;
  assign n4213 = n2343 | n3715 ;
  assign n4214 = n394 | n4213 ;
  assign n4215 = n972 | n4214 ;
  assign n4216 = n2197 | n4215 ;
  assign n4217 = n1525 | n4216 ;
  assign n4218 = n751 | n4217 ;
  assign n4219 = n352 | n4218 ;
  assign n4220 = n314 | n4219 ;
  assign n4221 = n172 | n4220 ;
  assign n4222 = n367 | n4221 ;
  assign n4223 = n108 | n4222 ;
  assign n4224 = n256 | n4223 ;
  assign n4225 = n236 | n4224 ;
  assign n6467 = ~n4120 ;
  assign n4122 = n287 & n6467 ;
  assign n4229 = n5502 & n4120 ;
  assign n4230 = n4122 | n4229 ;
  assign n4232 = n4190 & n4230 ;
  assign n4226 = n3902 | n4041 ;
  assign n4227 = n4040 & n4226 ;
  assign n4228 = n4039 | n4227 ;
  assign n4233 = n4193 & n4228 ;
  assign n4234 = n4232 | n4233 ;
  assign n4235 = n4175 & n4184 ;
  assign n4236 = n4127 & n4187 ;
  assign n4237 = n4235 | n4236 ;
  assign n3951 = n3324 & n6409 ;
  assign n6468 = ~n4109 ;
  assign n4110 = n3248 & n6468 ;
  assign n4238 = n3951 | n4110 ;
  assign n4239 = n287 | n4238 ;
  assign n4240 = n287 & n4238 ;
  assign n6469 = ~n4240 ;
  assign n4241 = n4239 & n6469 ;
  assign n3398 = n2891 & n6283 ;
  assign n2878 = n2558 & n2870 ;
  assign n3338 = n2879 & n3335 ;
  assign n4242 = n2878 | n3338 ;
  assign n4243 = n2860 & n6272 ;
  assign n4244 = n4242 | n4243 ;
  assign n4245 = n3398 | n4244 ;
  assign n6470 = ~n4245 ;
  assign n4246 = n1052 & n6470 ;
  assign n4247 = n5595 & n4245 ;
  assign n4248 = n4246 | n4247 ;
  assign n4249 = n4153 & n4162 ;
  assign n4250 = n4137 & n4165 ;
  assign n4251 = n4249 | n4250 ;
  assign n4252 = n4141 & n4150 ;
  assign n6471 = ~n4146 ;
  assign n4253 = n523 & n6471 ;
  assign n4254 = n2611 & n4253 ;
  assign n4255 = n4252 | n4254 ;
  assign n2609 = n523 & n6109 ;
  assign n2697 = n6091 & n2693 ;
  assign n2834 = n2598 & n2831 ;
  assign n4256 = n2697 | n2834 ;
  assign n4257 = n2589 & n2699 ;
  assign n4258 = n4256 | n4257 ;
  assign n4259 = n2713 & n6165 ;
  assign n4260 = n4258 | n4259 ;
  assign n4261 = n2609 | n4260 ;
  assign n4262 = n2609 & n4260 ;
  assign n6472 = ~n4262 ;
  assign n4263 = n4261 & n6472 ;
  assign n4264 = n4255 & n4263 ;
  assign n4265 = n4255 | n4263 ;
  assign n6473 = ~n4264 ;
  assign n4266 = n6473 & n4265 ;
  assign n2750 = n6081 & n2748 ;
  assign n4267 = n2584 & n2733 ;
  assign n4268 = n2564 & n2742 ;
  assign n4269 = n4267 | n4268 ;
  assign n4270 = n2750 | n4269 ;
  assign n4271 = n2727 & n6213 ;
  assign n4272 = n4270 | n4271 ;
  assign n4273 = n672 & n4272 ;
  assign n4274 = n672 | n4272 ;
  assign n6474 = ~n4273 ;
  assign n4275 = n6474 & n4274 ;
  assign n6475 = ~n4266 ;
  assign n4276 = n6475 & n4275 ;
  assign n6476 = ~n4275 ;
  assign n4277 = n4266 & n6476 ;
  assign n4278 = n4276 | n4277 ;
  assign n6477 = ~n4251 ;
  assign n4279 = n6477 & n4278 ;
  assign n6478 = ~n4278 ;
  assign n4281 = n4251 & n6478 ;
  assign n4282 = n4279 | n4281 ;
  assign n6479 = ~n4248 ;
  assign n4283 = n6479 & n4282 ;
  assign n6480 = ~n4282 ;
  assign n4284 = n4248 & n6480 ;
  assign n4285 = n4283 | n4284 ;
  assign n4286 = n4170 | n4174 ;
  assign n4287 = n4285 | n4286 ;
  assign n4288 = n4285 & n4286 ;
  assign n6481 = ~n4288 ;
  assign n4289 = n4287 & n6481 ;
  assign n3808 = n292 & n6372 ;
  assign n4290 = n2562 & n3314 ;
  assign n4291 = n2574 & n3673 ;
  assign n4292 = n4290 | n4291 ;
  assign n4293 = n3808 | n4292 ;
  assign n4294 = n2581 | n4293 ;
  assign n6482 = ~n4293 ;
  assign n4295 = n3824 & n6482 ;
  assign n6483 = ~n4295 ;
  assign n4296 = n4294 & n6483 ;
  assign n4297 = n274 & n4296 ;
  assign n4298 = n274 | n4296 ;
  assign n6484 = ~n4297 ;
  assign n4299 = n6484 & n4298 ;
  assign n4300 = n4289 & n4299 ;
  assign n4301 = n4289 | n4299 ;
  assign n6485 = ~n4300 ;
  assign n4302 = n6485 & n4301 ;
  assign n4303 = n4241 & n4302 ;
  assign n4304 = n4241 | n4302 ;
  assign n6486 = ~n4303 ;
  assign n4305 = n6486 & n4304 ;
  assign n4306 = n4237 & n4305 ;
  assign n4307 = n4237 | n4305 ;
  assign n6487 = ~n4306 ;
  assign n4308 = n6487 & n4307 ;
  assign n4309 = n4234 & n4308 ;
  assign n4310 = n4234 | n4308 ;
  assign n6488 = ~n4309 ;
  assign n4311 = n6488 & n4310 ;
  assign n6489 = ~n4311 ;
  assign n4312 = n4225 & n6489 ;
  assign n6490 = ~n4225 ;
  assign n4313 = n6490 & n4311 ;
  assign n4314 = n4312 | n4313 ;
  assign n4315 = n4202 & n4314 ;
  assign n4316 = n4202 | n4313 ;
  assign n4317 = n4312 | n4316 ;
  assign n6491 = ~n4315 ;
  assign n4318 = n6491 & n4317 ;
  assign n4319 = n4206 & n4318 ;
  assign n4320 = n4206 | n4318 ;
  assign n6492 = ~n4319 ;
  assign n4321 = n6492 & n4320 ;
  assign n4322 = n4207 | n4208 ;
  assign n4323 = n4077 & n4322 ;
  assign n4324 = n4321 & n4323 ;
  assign n4325 = n4321 | n4323 ;
  assign n6493 = ~n4324 ;
  assign n28 = n6493 & n4325 ;
  assign n4327 = n4225 & n4311 ;
  assign n4328 = n4315 | n4327 ;
  assign n4329 = n343 | n495 ;
  assign n4330 = n298 | n4329 ;
  assign n4331 = n2469 | n4330 ;
  assign n4332 = n1001 | n4331 ;
  assign n4333 = n768 | n4332 ;
  assign n4334 = n643 | n4333 ;
  assign n4335 = n2423 | n4334 ;
  assign n4336 = n175 | n4335 ;
  assign n4337 = n192 | n4336 ;
  assign n4338 = n588 | n4337 ;
  assign n4339 = n4306 | n4309 ;
  assign n4340 = n4300 | n4303 ;
  assign n4341 = n4248 & n4282 ;
  assign n4342 = n4288 | n4341 ;
  assign n4280 = n4251 & n4278 ;
  assign n4343 = n4266 & n4275 ;
  assign n4344 = n4280 | n4343 ;
  assign n2698 = n2589 & n2693 ;
  assign n2835 = n6091 & n2831 ;
  assign n4345 = n2698 | n2835 ;
  assign n4346 = n2584 & n2699 ;
  assign n4347 = n4345 | n4346 ;
  assign n4348 = n2713 & n3051 ;
  assign n4349 = n4347 | n4348 ;
  assign n6494 = ~n4349 ;
  assign n4350 = n523 & n6494 ;
  assign n4351 = n5542 & n4349 ;
  assign n4352 = n4350 | n4351 ;
  assign n4353 = n287 & n523 ;
  assign n4354 = n2598 & n4353 ;
  assign n6495 = ~n4354 ;
  assign n4355 = n287 & n6495 ;
  assign n6496 = ~n4353 ;
  assign n4356 = n2598 & n6496 ;
  assign n4357 = n523 & n4356 ;
  assign n4358 = n4355 | n4357 ;
  assign n4359 = n4352 | n4358 ;
  assign n4360 = n4352 & n4358 ;
  assign n6497 = ~n4360 ;
  assign n4361 = n4359 & n6497 ;
  assign n4362 = n523 & n2605 ;
  assign n6498 = ~n4260 ;
  assign n4363 = n6498 & n4362 ;
  assign n4364 = n4264 | n4363 ;
  assign n4365 = n4361 | n4364 ;
  assign n4366 = n4361 & n4364 ;
  assign n6499 = ~n4366 ;
  assign n4367 = n4365 & n6499 ;
  assign n2729 = n6124 & n2727 ;
  assign n2738 = n2564 & n2733 ;
  assign n2746 = n6081 & n2742 ;
  assign n4368 = n2738 | n2746 ;
  assign n4369 = n2558 & n2748 ;
  assign n4370 = n4368 | n4369 ;
  assign n4371 = n2729 | n4370 ;
  assign n6500 = ~n4371 ;
  assign n4372 = n672 & n6500 ;
  assign n4373 = n5514 & n4371 ;
  assign n4374 = n4372 | n4373 ;
  assign n6501 = ~n4367 ;
  assign n4375 = n6501 & n4374 ;
  assign n6502 = ~n4374 ;
  assign n4376 = n4367 & n6502 ;
  assign n4377 = n4375 | n4376 ;
  assign n4378 = n4344 | n4377 ;
  assign n4379 = n4344 & n4377 ;
  assign n6503 = ~n4379 ;
  assign n4380 = n4378 & n6503 ;
  assign n3381 = n2891 & n6278 ;
  assign n3339 = n2870 & n3335 ;
  assign n3349 = n2879 & n6272 ;
  assign n4381 = n3339 | n3349 ;
  assign n4382 = n2860 & n3314 ;
  assign n4383 = n4381 | n4382 ;
  assign n4384 = n3381 | n4383 ;
  assign n6504 = ~n4384 ;
  assign n4385 = n1052 & n6504 ;
  assign n4386 = n5595 & n4384 ;
  assign n4387 = n4385 | n4386 ;
  assign n4388 = n4380 | n4387 ;
  assign n4389 = n4380 & n4387 ;
  assign n6505 = ~n4389 ;
  assign n4390 = n4388 & n6505 ;
  assign n6506 = ~n4342 ;
  assign n4391 = n6506 & n4390 ;
  assign n6507 = ~n4390 ;
  assign n4392 = n4342 & n6507 ;
  assign n4393 = n4391 | n4392 ;
  assign n3967 = n2581 & n3965 ;
  assign n3678 = n2562 & n3673 ;
  assign n3811 = n2574 & n6372 ;
  assign n4394 = n3678 | n3811 ;
  assign n4395 = n292 & n6409 ;
  assign n4396 = n4394 | n4395 ;
  assign n4397 = n3967 | n4396 ;
  assign n6508 = ~n4397 ;
  assign n4398 = n274 & n6508 ;
  assign n4399 = n5721 & n4397 ;
  assign n4400 = n4398 | n4399 ;
  assign n4401 = n4393 & n4400 ;
  assign n4402 = n4393 | n4400 ;
  assign n6509 = ~n4401 ;
  assign n4403 = n6509 & n4402 ;
  assign n4404 = n4340 & n4403 ;
  assign n4405 = n4340 | n4403 ;
  assign n6510 = ~n4404 ;
  assign n4406 = n6510 & n4405 ;
  assign n6511 = ~n4339 ;
  assign n4407 = n6511 & n4406 ;
  assign n6512 = ~n4406 ;
  assign n4408 = n4339 & n6512 ;
  assign n4409 = n4407 | n4408 ;
  assign n6513 = ~n4338 ;
  assign n4410 = n6513 & n4409 ;
  assign n6514 = ~n4409 ;
  assign n4411 = n4338 & n6514 ;
  assign n4412 = n4410 | n4411 ;
  assign n4413 = n4328 | n4412 ;
  assign n4414 = n4328 & n4412 ;
  assign n6515 = ~n4414 ;
  assign n4415 = n4413 & n6515 ;
  assign n4416 = n4319 & n4415 ;
  assign n4417 = n4319 | n4415 ;
  assign n6516 = ~n4416 ;
  assign n4418 = n6516 & n4417 ;
  assign n4419 = n4321 | n4322 ;
  assign n4420 = n4077 & n4419 ;
  assign n4421 = n4418 & n4420 ;
  assign n4422 = n4418 | n4420 ;
  assign n6517 = ~n4421 ;
  assign n29 = n6517 & n4422 ;
  assign n4424 = n4338 & n4409 ;
  assign n4425 = n4414 | n4424 ;
  assign n4426 = n314 | n356 ;
  assign n4427 = n471 | n4426 ;
  assign n4428 = n187 | n823 ;
  assign n4429 = n4427 | n4428 ;
  assign n4430 = n2320 | n4429 ;
  assign n4431 = n311 | n4430 ;
  assign n4432 = n3934 | n4431 ;
  assign n4433 = n3285 | n4432 ;
  assign n4434 = n4053 | n4433 ;
  assign n4435 = n366 | n4434 ;
  assign n4436 = n175 | n4435 ;
  assign n4437 = n414 | n4436 ;
  assign n4438 = n296 | n4437 ;
  assign n4439 = n235 | n4438 ;
  assign n4440 = n4124 & n4190 ;
  assign n4231 = n4190 | n4230 ;
  assign n6518 = ~n4232 ;
  assign n4441 = n4231 & n6518 ;
  assign n4442 = n4103 & n4441 ;
  assign n4443 = n4440 | n4442 ;
  assign n4444 = n4307 & n4443 ;
  assign n4445 = n4306 | n4444 ;
  assign n4446 = n4406 & n4445 ;
  assign n4447 = n4404 | n4446 ;
  assign n4448 = n4342 & n4390 ;
  assign n4449 = n4401 | n4448 ;
  assign n4117 = n2581 & n4115 ;
  assign n4501 = n2562 & n6372 ;
  assign n4502 = n2574 & n6409 ;
  assign n4503 = n4501 | n4502 ;
  assign n4504 = n4117 | n4503 ;
  assign n6519 = ~n4504 ;
  assign n4505 = n274 & n6519 ;
  assign n4506 = n5721 & n4504 ;
  assign n4507 = n4505 | n4506 ;
  assign n4450 = n4379 | n4389 ;
  assign n3697 = n2891 & n3696 ;
  assign n3321 = n2879 & n3314 ;
  assign n3350 = n2870 & n6272 ;
  assign n4486 = n3321 | n3350 ;
  assign n4487 = n2860 & n3673 ;
  assign n4488 = n4486 | n4487 ;
  assign n4489 = n3697 | n4488 ;
  assign n4490 = n1052 | n4489 ;
  assign n4491 = n1052 & n4489 ;
  assign n6520 = ~n4491 ;
  assign n4492 = n4490 & n6520 ;
  assign n4451 = n4367 & n4374 ;
  assign n4452 = n4366 | n4451 ;
  assign n3416 = n2727 & n3412 ;
  assign n2734 = n6081 & n2733 ;
  assign n2747 = n2558 & n2742 ;
  assign n4473 = n2734 | n2747 ;
  assign n4474 = n2748 & n3335 ;
  assign n4475 = n4473 | n4474 ;
  assign n4476 = n3416 | n4475 ;
  assign n6521 = ~n4476 ;
  assign n4477 = n672 & n6521 ;
  assign n4478 = n5514 & n4476 ;
  assign n4479 = n4477 | n4478 ;
  assign n4453 = n4354 | n4360 ;
  assign n4454 = n6091 & n4353 ;
  assign n6522 = ~n4454 ;
  assign n4455 = n287 & n6522 ;
  assign n4456 = n2594 | n4353 ;
  assign n6523 = ~n4456 ;
  assign n4457 = n523 & n6523 ;
  assign n4458 = n4455 | n4457 ;
  assign n4459 = n4453 | n4458 ;
  assign n4460 = n4453 & n4458 ;
  assign n6524 = ~n4460 ;
  assign n4461 = n4459 & n6524 ;
  assign n2705 = n2564 & n2699 ;
  assign n4462 = n2584 & n2693 ;
  assign n4463 = n2589 & n2831 ;
  assign n4464 = n4462 | n4463 ;
  assign n4465 = n2705 | n4464 ;
  assign n4466 = n2713 & n3093 ;
  assign n4467 = n4465 | n4466 ;
  assign n4468 = n523 & n4467 ;
  assign n4469 = n523 | n4467 ;
  assign n6525 = ~n4468 ;
  assign n4470 = n6525 & n4469 ;
  assign n6526 = ~n4461 ;
  assign n4471 = n6526 & n4470 ;
  assign n6527 = ~n4470 ;
  assign n4472 = n4461 & n6527 ;
  assign n4480 = n4471 | n4472 ;
  assign n4481 = n4479 & n4480 ;
  assign n4482 = n4471 | n4479 ;
  assign n4483 = n4472 | n4482 ;
  assign n6528 = ~n4481 ;
  assign n4484 = n6528 & n4483 ;
  assign n6529 = ~n4484 ;
  assign n4485 = n4452 & n6529 ;
  assign n6530 = ~n4452 ;
  assign n4493 = n6530 & n4484 ;
  assign n4494 = n4485 | n4493 ;
  assign n4495 = n4492 & n4494 ;
  assign n4496 = n4492 | n4493 ;
  assign n4497 = n4485 | n4496 ;
  assign n6531 = ~n4495 ;
  assign n4498 = n6531 & n4497 ;
  assign n6532 = ~n4498 ;
  assign n4499 = n4450 & n6532 ;
  assign n6533 = ~n4450 ;
  assign n4500 = n6533 & n4498 ;
  assign n4508 = n4499 | n4500 ;
  assign n4509 = n4507 & n4508 ;
  assign n4510 = n4500 | n4507 ;
  assign n4511 = n4499 | n4510 ;
  assign n6534 = ~n4509 ;
  assign n4512 = n6534 & n4511 ;
  assign n4513 = n4449 & n4512 ;
  assign n4514 = n4449 | n4512 ;
  assign n6535 = ~n4513 ;
  assign n4515 = n6535 & n4514 ;
  assign n6536 = ~n4447 ;
  assign n4516 = n6536 & n4515 ;
  assign n6537 = ~n4515 ;
  assign n4517 = n4447 & n6537 ;
  assign n4518 = n4516 | n4517 ;
  assign n4519 = n4439 | n4518 ;
  assign n4520 = n4439 & n4518 ;
  assign n6538 = ~n4520 ;
  assign n4521 = n4519 & n6538 ;
  assign n6539 = ~n4425 ;
  assign n4522 = n6539 & n4521 ;
  assign n6540 = ~n4521 ;
  assign n4523 = n4425 & n6540 ;
  assign n4524 = n4522 | n4523 ;
  assign n4525 = n4416 & n4524 ;
  assign n4526 = n4416 | n4524 ;
  assign n6541 = ~n4525 ;
  assign n4527 = n6541 & n4526 ;
  assign n4528 = n4418 | n4419 ;
  assign n4529 = n4077 & n4528 ;
  assign n4530 = n4527 & n4529 ;
  assign n4531 = n4527 | n4529 ;
  assign n6542 = ~n4530 ;
  assign n30 = n6542 & n4531 ;
  assign n4533 = n4425 & n4521 ;
  assign n4534 = n4520 | n4533 ;
  assign n4535 = n313 | n1164 ;
  assign n4536 = n585 | n4535 ;
  assign n4537 = n2426 | n4536 ;
  assign n4538 = n2343 | n4537 ;
  assign n4539 = n153 | n4538 ;
  assign n4540 = n366 | n4539 ;
  assign n4541 = n1002 | n4540 ;
  assign n4542 = n354 | n4541 ;
  assign n4543 = n251 | n996 ;
  assign n4544 = n2463 | n4543 ;
  assign n4545 = n3301 | n4544 ;
  assign n4546 = n4542 | n4545 ;
  assign n4547 = n334 | n4546 ;
  assign n4548 = n147 | n4547 ;
  assign n4549 = n169 | n4548 ;
  assign n4550 = n166 | n4549 ;
  assign n4551 = n446 | n4550 ;
  assign n4552 = n145 | n4551 ;
  assign n4553 = n4339 & n4405 ;
  assign n4554 = n4404 | n4553 ;
  assign n4555 = n4515 & n4554 ;
  assign n4556 = n4513 | n4555 ;
  assign n4557 = n4450 & n4498 ;
  assign n4558 = n4509 | n4557 ;
  assign n4559 = n4452 & n4484 ;
  assign n4560 = n4495 | n4559 ;
  assign n3948 = n2562 & n6409 ;
  assign n4111 = n2581 & n6468 ;
  assign n4561 = n3948 | n4111 ;
  assign n6543 = ~n4561 ;
  assign n4562 = n274 & n6543 ;
  assign n4563 = n5721 & n4561 ;
  assign n4564 = n4562 | n4563 ;
  assign n4565 = n4560 | n4564 ;
  assign n4566 = n4560 & n4564 ;
  assign n6544 = ~n4566 ;
  assign n4567 = n4565 & n6544 ;
  assign n3826 = n2891 & n6375 ;
  assign n3318 = n2870 & n3314 ;
  assign n3679 = n2879 & n3673 ;
  assign n4568 = n3318 | n3679 ;
  assign n4569 = n2860 & n6372 ;
  assign n4570 = n4568 | n4569 ;
  assign n4571 = n3826 | n4570 ;
  assign n6545 = ~n4571 ;
  assign n4572 = n1052 & n6545 ;
  assign n4573 = n5595 & n4571 ;
  assign n4574 = n4572 | n4573 ;
  assign n4575 = n4461 & n4470 ;
  assign n4576 = n4481 | n4575 ;
  assign n3397 = n2727 & n6283 ;
  assign n2741 = n2558 & n2733 ;
  assign n3340 = n2742 & n3335 ;
  assign n4597 = n2741 | n3340 ;
  assign n4598 = n2748 & n6272 ;
  assign n4599 = n4597 | n4598 ;
  assign n4600 = n3397 | n4599 ;
  assign n6546 = ~n4600 ;
  assign n4601 = n672 & n6546 ;
  assign n4602 = n5514 & n4600 ;
  assign n4603 = n4601 | n4602 ;
  assign n4577 = n4454 | n4460 ;
  assign n4578 = n2589 & n4353 ;
  assign n6547 = ~n4578 ;
  assign n4579 = n287 & n6547 ;
  assign n4580 = n2589 & n6496 ;
  assign n4581 = n523 & n4580 ;
  assign n4582 = n4579 | n4581 ;
  assign n4583 = n4577 | n4582 ;
  assign n4584 = n4577 & n4582 ;
  assign n6548 = ~n4584 ;
  assign n4585 = n4583 & n6548 ;
  assign n2706 = n6081 & n2699 ;
  assign n4586 = n2564 & n2693 ;
  assign n4587 = n2584 & n2831 ;
  assign n4588 = n4586 | n4587 ;
  assign n4589 = n2706 | n4588 ;
  assign n4590 = n2713 & n6213 ;
  assign n4591 = n4589 | n4590 ;
  assign n4592 = n523 & n4591 ;
  assign n4593 = n523 | n4591 ;
  assign n6549 = ~n4592 ;
  assign n4594 = n6549 & n4593 ;
  assign n6550 = ~n4585 ;
  assign n4595 = n6550 & n4594 ;
  assign n6551 = ~n4594 ;
  assign n4596 = n4585 & n6551 ;
  assign n4604 = n4595 | n4596 ;
  assign n4605 = n4603 & n4604 ;
  assign n4606 = n4595 | n4603 ;
  assign n4607 = n4596 | n4606 ;
  assign n6552 = ~n4605 ;
  assign n4608 = n6552 & n4607 ;
  assign n6553 = ~n4608 ;
  assign n4609 = n4576 & n6553 ;
  assign n6554 = ~n4576 ;
  assign n4610 = n6554 & n4608 ;
  assign n4611 = n4609 | n4610 ;
  assign n4612 = n4574 & n4611 ;
  assign n4613 = n4574 | n4610 ;
  assign n4614 = n4609 | n4613 ;
  assign n6555 = ~n4612 ;
  assign n4615 = n6555 & n4614 ;
  assign n6556 = ~n4567 ;
  assign n4616 = n6556 & n4615 ;
  assign n6557 = ~n4615 ;
  assign n4617 = n4567 & n6557 ;
  assign n4618 = n4616 | n4617 ;
  assign n4619 = n4558 & n4618 ;
  assign n4620 = n4558 | n4618 ;
  assign n6558 = ~n4619 ;
  assign n4621 = n6558 & n4620 ;
  assign n6559 = ~n4556 ;
  assign n4622 = n6559 & n4621 ;
  assign n6560 = ~n4621 ;
  assign n4623 = n4556 & n6560 ;
  assign n4624 = n4622 | n4623 ;
  assign n6561 = ~n4552 ;
  assign n4625 = n6561 & n4624 ;
  assign n6562 = ~n4624 ;
  assign n4626 = n4552 & n6562 ;
  assign n4627 = n4625 | n4626 ;
  assign n4628 = n4534 | n4627 ;
  assign n4629 = n4534 & n4627 ;
  assign n6563 = ~n4629 ;
  assign n4630 = n4628 & n6563 ;
  assign n4631 = n4525 & n4630 ;
  assign n4632 = n4525 | n4630 ;
  assign n6564 = ~n4631 ;
  assign n4633 = n6564 & n4632 ;
  assign n4634 = n4527 | n4528 ;
  assign n4635 = n4077 & n4634 ;
  assign n4636 = n4633 & n4635 ;
  assign n4637 = n4633 | n4635 ;
  assign n6565 = ~n4636 ;
  assign n31 = n6565 & n4637 ;
  assign n4639 = n4552 & n4624 ;
  assign n4640 = n4629 | n4639 ;
  assign n4641 = n4567 & n4615 ;
  assign n4642 = n4566 | n4641 ;
  assign n4643 = n4576 & n4608 ;
  assign n4644 = n4612 | n4643 ;
  assign n3953 = n2860 & n6409 ;
  assign n4645 = n2870 & n3673 ;
  assign n4646 = n2879 & n6372 ;
  assign n4647 = n4645 | n4646 ;
  assign n4648 = n3953 | n4647 ;
  assign n4649 = n2891 & n3965 ;
  assign n4650 = n4648 | n4649 ;
  assign n4651 = n1052 & n4650 ;
  assign n4652 = n1052 | n4650 ;
  assign n6566 = ~n4651 ;
  assign n4653 = n6566 & n4652 ;
  assign n4654 = n4644 & n4653 ;
  assign n4655 = n4644 | n4653 ;
  assign n6567 = ~n4654 ;
  assign n4656 = n6567 & n4655 ;
  assign n4657 = n4585 & n4594 ;
  assign n4658 = n4605 | n4657 ;
  assign n4659 = n4578 | n4584 ;
  assign n2714 = n6124 & n2713 ;
  assign n2696 = n6081 & n2693 ;
  assign n2836 = n2564 & n2831 ;
  assign n4660 = n2696 | n2836 ;
  assign n4661 = n2558 & n2699 ;
  assign n4662 = n4660 | n4661 ;
  assign n4663 = n2714 | n4662 ;
  assign n6568 = ~n4663 ;
  assign n4664 = n523 & n6568 ;
  assign n4665 = n5542 & n4663 ;
  assign n4666 = n4664 | n4665 ;
  assign n4667 = n523 & n2584 ;
  assign n289 = n274 | n287 ;
  assign n4668 = n274 & n287 ;
  assign n6569 = ~n4668 ;
  assign n4669 = n289 & n6569 ;
  assign n4670 = n4667 & n4669 ;
  assign n4671 = n4667 | n4669 ;
  assign n6570 = ~n4670 ;
  assign n4672 = n6570 & n4671 ;
  assign n6571 = ~n4666 ;
  assign n4673 = n6571 & n4672 ;
  assign n6572 = ~n4672 ;
  assign n4674 = n4666 & n6572 ;
  assign n4675 = n4673 | n4674 ;
  assign n4676 = n4659 | n4675 ;
  assign n4677 = n4659 & n4675 ;
  assign n6573 = ~n4677 ;
  assign n4678 = n4676 & n6573 ;
  assign n3316 = n2748 & n3314 ;
  assign n4679 = n2733 & n3335 ;
  assign n4680 = n2742 & n6272 ;
  assign n4681 = n4679 | n4680 ;
  assign n4682 = n3316 | n4681 ;
  assign n4683 = n2727 & n6278 ;
  assign n4684 = n4682 | n4683 ;
  assign n4685 = n672 & n4684 ;
  assign n4686 = n672 | n4684 ;
  assign n6574 = ~n4685 ;
  assign n4687 = n6574 & n4686 ;
  assign n6575 = ~n4678 ;
  assign n4688 = n6575 & n4687 ;
  assign n6576 = ~n4687 ;
  assign n4689 = n4678 & n6576 ;
  assign n4690 = n4688 | n4689 ;
  assign n6577 = ~n4690 ;
  assign n4691 = n4658 & n6577 ;
  assign n6578 = ~n4658 ;
  assign n4692 = n6578 & n4690 ;
  assign n4693 = n4691 | n4692 ;
  assign n6579 = ~n4693 ;
  assign n4694 = n4656 & n6579 ;
  assign n6580 = ~n4656 ;
  assign n4695 = n6580 & n4693 ;
  assign n4696 = n4694 | n4695 ;
  assign n4697 = n4642 | n4696 ;
  assign n4698 = n4642 & n4696 ;
  assign n6581 = ~n4698 ;
  assign n4699 = n4697 & n6581 ;
  assign n4700 = n4447 & n4514 ;
  assign n4701 = n4513 | n4700 ;
  assign n4702 = n4621 & n4701 ;
  assign n4703 = n4619 | n4702 ;
  assign n6582 = ~n4703 ;
  assign n4704 = n4699 & n6582 ;
  assign n6583 = ~n4699 ;
  assign n4705 = n6583 & n4703 ;
  assign n4706 = n4704 | n4705 ;
  assign n4707 = n957 | n2283 ;
  assign n4708 = n4427 | n4707 ;
  assign n4709 = n825 | n4708 ;
  assign n4710 = n4542 | n4709 ;
  assign n4711 = n126 | n4710 ;
  assign n4712 = n192 | n4711 ;
  assign n4713 = n134 | n4712 ;
  assign n4714 = n216 | n4713 ;
  assign n4715 = n1137 | n4714 ;
  assign n4716 = n165 | n4715 ;
  assign n4717 = n444 | n4716 ;
  assign n4718 = n4706 | n4717 ;
  assign n4719 = n4706 & n4717 ;
  assign n6584 = ~n4719 ;
  assign n4720 = n4718 & n6584 ;
  assign n6585 = ~n4640 ;
  assign n4721 = n6585 & n4720 ;
  assign n6586 = ~n4720 ;
  assign n4722 = n4640 & n6586 ;
  assign n4723 = n4721 | n4722 ;
  assign n4724 = n4631 & n4723 ;
  assign n4725 = n4631 | n4723 ;
  assign n6587 = ~n4724 ;
  assign n4726 = n6587 & n4725 ;
  assign n4727 = n4633 | n4634 ;
  assign n4728 = n4077 & n4727 ;
  assign n4729 = n4726 & n4728 ;
  assign n4730 = n4726 | n4728 ;
  assign n6588 = ~n4729 ;
  assign n32 = n6588 & n4730 ;
  assign n4732 = n4640 & n4720 ;
  assign n4733 = n4719 | n4732 ;
  assign n4734 = n608 | n2182 ;
  assign n4735 = n162 | n4734 ;
  assign n4736 = n219 | n4735 ;
  assign n4737 = n217 | n4736 ;
  assign n4738 = n164 | n4737 ;
  assign n4739 = n223 | n4738 ;
  assign n4740 = n445 | n4739 ;
  assign n4741 = n108 | n4740 ;
  assign n4742 = n209 | n4741 ;
  assign n4743 = n987 | n2345 ;
  assign n4744 = n1005 | n4743 ;
  assign n4745 = n3736 | n4744 ;
  assign n4746 = n4742 | n4745 ;
  assign n4747 = n405 | n4746 ;
  assign n4748 = n255 | n4747 ;
  assign n4749 = n205 | n4748 ;
  assign n4750 = n358 | n4749 ;
  assign n4751 = n222 | n4750 ;
  assign n4752 = n323 | n4751 ;
  assign n4753 = n468 | n4752 ;
  assign n4754 = n4699 & n4703 ;
  assign n4755 = n4698 | n4754 ;
  assign n4756 = n4656 & n4693 ;
  assign n4757 = n4654 | n4756 ;
  assign n4118 = n2891 & n4115 ;
  assign n4758 = n2870 & n6372 ;
  assign n4759 = n2879 & n6409 ;
  assign n4760 = n4758 | n4759 ;
  assign n4761 = n4118 | n4760 ;
  assign n6589 = ~n4761 ;
  assign n4762 = n1052 & n6589 ;
  assign n4763 = n5595 & n4761 ;
  assign n4764 = n4762 | n4763 ;
  assign n4765 = n4678 & n4687 ;
  assign n4766 = n4658 & n4690 ;
  assign n4767 = n4765 | n4766 ;
  assign n4768 = n4666 & n4672 ;
  assign n4769 = n4677 | n4768 ;
  assign n2567 = n523 & n2564 ;
  assign n4770 = n289 & n6570 ;
  assign n4771 = n2567 & n4770 ;
  assign n4772 = n2567 | n4770 ;
  assign n6590 = ~n4771 ;
  assign n4773 = n6590 & n4772 ;
  assign n3337 = n2699 & n3335 ;
  assign n4774 = n2558 & n2693 ;
  assign n4775 = n6081 & n2831 ;
  assign n4776 = n4774 | n4775 ;
  assign n4777 = n3337 | n4776 ;
  assign n4778 = n2713 & n3412 ;
  assign n4779 = n4777 | n4778 ;
  assign n4780 = n523 & n4779 ;
  assign n4781 = n523 | n4779 ;
  assign n6591 = ~n4780 ;
  assign n4782 = n6591 & n4781 ;
  assign n6592 = ~n4773 ;
  assign n4783 = n6592 & n4782 ;
  assign n6593 = ~n4782 ;
  assign n4785 = n4773 & n6593 ;
  assign n4786 = n4783 | n4785 ;
  assign n6594 = ~n4786 ;
  assign n4788 = n4769 & n6594 ;
  assign n6595 = ~n4769 ;
  assign n4789 = n6595 & n4786 ;
  assign n4790 = n4788 | n4789 ;
  assign n3698 = n2727 & n3696 ;
  assign n3315 = n2742 & n3314 ;
  assign n3351 = n2733 & n6272 ;
  assign n4791 = n3315 | n3351 ;
  assign n4792 = n2748 & n3673 ;
  assign n4793 = n4791 | n4792 ;
  assign n4794 = n3698 | n4793 ;
  assign n6596 = ~n4794 ;
  assign n4795 = n672 & n6596 ;
  assign n4796 = n5514 & n4794 ;
  assign n4797 = n4795 | n4796 ;
  assign n4798 = n4790 & n4797 ;
  assign n4799 = n4789 | n4797 ;
  assign n4800 = n4788 | n4799 ;
  assign n6597 = ~n4798 ;
  assign n4801 = n6597 & n4800 ;
  assign n6598 = ~n4767 ;
  assign n4802 = n6598 & n4801 ;
  assign n6599 = ~n4801 ;
  assign n4803 = n4767 & n6599 ;
  assign n4804 = n4802 | n4803 ;
  assign n6600 = ~n4764 ;
  assign n4805 = n6600 & n4804 ;
  assign n6601 = ~n4804 ;
  assign n4806 = n4764 & n6601 ;
  assign n4807 = n4805 | n4806 ;
  assign n4808 = n4757 & n4807 ;
  assign n4809 = n4757 | n4807 ;
  assign n6602 = ~n4808 ;
  assign n4810 = n6602 & n4809 ;
  assign n4811 = n4755 & n4810 ;
  assign n4812 = n4755 | n4810 ;
  assign n6603 = ~n4811 ;
  assign n4813 = n6603 & n4812 ;
  assign n6604 = ~n4753 ;
  assign n4814 = n6604 & n4813 ;
  assign n6605 = ~n4813 ;
  assign n4815 = n4753 & n6605 ;
  assign n4816 = n4814 | n4815 ;
  assign n6606 = ~n4816 ;
  assign n4817 = n4733 & n6606 ;
  assign n6607 = ~n4733 ;
  assign n4818 = n6607 & n4816 ;
  assign n4819 = n4817 | n4818 ;
  assign n4820 = n4724 & n4819 ;
  assign n4821 = n4724 | n4819 ;
  assign n6608 = ~n4820 ;
  assign n4822 = n6608 & n4821 ;
  assign n4823 = n4726 | n4727 ;
  assign n4824 = n4077 & n4823 ;
  assign n4825 = n4822 & n4824 ;
  assign n4826 = n4822 | n4824 ;
  assign n6609 = ~n4825 ;
  assign n33 = n6609 & n4826 ;
  assign n4828 = n4753 & n4813 ;
  assign n4829 = n4733 & n4816 ;
  assign n4830 = n4828 | n4829 ;
  assign n4831 = n773 | n825 ;
  assign n4832 = n202 | n4831 ;
  assign n4833 = n3273 | n4832 ;
  assign n4834 = n2437 | n4833 ;
  assign n4835 = n3301 | n4834 ;
  assign n4836 = n334 | n4835 ;
  assign n4837 = n324 | n4836 ;
  assign n4838 = n223 | n4837 ;
  assign n4839 = n130 | n4838 ;
  assign n4840 = n232 | n4839 ;
  assign n4841 = n353 | n4840 ;
  assign n4842 = n214 | n4841 ;
  assign n4843 = n4767 & n4801 ;
  assign n4844 = n4764 & n4804 ;
  assign n4845 = n4843 | n4844 ;
  assign n4784 = n4773 & n4782 ;
  assign n6610 = ~n4784 ;
  assign n4846 = n4772 & n6610 ;
  assign n3399 = n2713 & n6283 ;
  assign n2837 = n2558 & n2831 ;
  assign n3341 = n2693 & n3335 ;
  assign n4847 = n2837 | n3341 ;
  assign n4848 = n2699 & n6272 ;
  assign n4849 = n4847 | n4848 ;
  assign n4850 = n3399 | n4849 ;
  assign n6611 = ~n4850 ;
  assign n4851 = n523 & n6611 ;
  assign n4852 = n5542 & n4850 ;
  assign n4853 = n4851 | n4852 ;
  assign n4854 = n523 & n6120 ;
  assign n4855 = n4853 & n4854 ;
  assign n4856 = n4853 | n4854 ;
  assign n6612 = ~n4855 ;
  assign n4857 = n6612 & n4856 ;
  assign n4858 = n4846 & n4857 ;
  assign n4859 = n4846 | n4857 ;
  assign n6613 = ~n4858 ;
  assign n4860 = n6613 & n4859 ;
  assign n3827 = n2727 & n6375 ;
  assign n3323 = n2733 & n3314 ;
  assign n3680 = n2742 & n3673 ;
  assign n4861 = n3323 | n3680 ;
  assign n4862 = n2748 & n6372 ;
  assign n4863 = n4861 | n4862 ;
  assign n4864 = n3827 | n4863 ;
  assign n6614 = ~n4864 ;
  assign n4865 = n672 & n6614 ;
  assign n4866 = n5514 & n4864 ;
  assign n4867 = n4865 | n4866 ;
  assign n6615 = ~n4860 ;
  assign n4868 = n6615 & n4867 ;
  assign n6616 = ~n4867 ;
  assign n4869 = n4860 & n6616 ;
  assign n4870 = n4868 | n4869 ;
  assign n4787 = n4769 & n4786 ;
  assign n4871 = n4787 | n4798 ;
  assign n3952 = n2870 & n6409 ;
  assign n4112 = n2891 & n6468 ;
  assign n4872 = n3952 | n4112 ;
  assign n6617 = ~n4872 ;
  assign n4873 = n1052 & n6617 ;
  assign n4874 = n5595 & n4872 ;
  assign n4875 = n4873 | n4874 ;
  assign n4876 = n4871 | n4875 ;
  assign n4877 = n4871 & n4875 ;
  assign n6618 = ~n4877 ;
  assign n4878 = n4876 & n6618 ;
  assign n6619 = ~n4870 ;
  assign n4879 = n6619 & n4878 ;
  assign n6620 = ~n4878 ;
  assign n4880 = n4870 & n6620 ;
  assign n4881 = n4879 | n4880 ;
  assign n4882 = n4845 | n4881 ;
  assign n4883 = n4845 & n4881 ;
  assign n6621 = ~n4883 ;
  assign n4884 = n4882 & n6621 ;
  assign n4885 = n4808 | n4811 ;
  assign n6622 = ~n4885 ;
  assign n4886 = n4884 & n6622 ;
  assign n6623 = ~n4884 ;
  assign n4887 = n6623 & n4885 ;
  assign n4888 = n4886 | n4887 ;
  assign n4889 = n4842 | n4888 ;
  assign n4890 = n4842 & n4888 ;
  assign n6624 = ~n4890 ;
  assign n4891 = n4889 & n6624 ;
  assign n6625 = ~n4830 ;
  assign n4892 = n6625 & n4891 ;
  assign n6626 = ~n4891 ;
  assign n4893 = n4830 & n6626 ;
  assign n4894 = n4892 | n4893 ;
  assign n4895 = n4820 & n4894 ;
  assign n4896 = n4820 | n4894 ;
  assign n6627 = ~n4895 ;
  assign n4897 = n6627 & n4896 ;
  assign n4898 = n4822 | n4823 ;
  assign n4899 = n4077 & n4898 ;
  assign n4900 = n4897 & n4899 ;
  assign n4901 = n4897 | n4899 ;
  assign n6628 = ~n4900 ;
  assign n34 = n6628 & n4901 ;
  assign n4903 = n4830 & n4891 ;
  assign n4904 = n4890 | n4903 ;
  assign n4905 = n257 | n654 ;
  assign n4906 = n475 | n4905 ;
  assign n4907 = n504 | n4906 ;
  assign n4908 = n208 | n4907 ;
  assign n4909 = n3724 | n4908 ;
  assign n4910 = n1151 | n4909 ;
  assign n4911 = n3301 | n4910 ;
  assign n4912 = n1003 | n4911 ;
  assign n4913 = n309 | n4912 ;
  assign n4914 = n190 | n4913 ;
  assign n4915 = n312 | n4914 ;
  assign n4916 = n4884 & n4885 ;
  assign n4917 = n4883 | n4916 ;
  assign n4918 = n4870 & n4878 ;
  assign n4919 = n4877 | n4918 ;
  assign n6629 = ~n4854 ;
  assign n4920 = n4853 & n6629 ;
  assign n4921 = n2567 | n2570 ;
  assign n6630 = ~n4921 ;
  assign n4922 = n523 & n6630 ;
  assign n4923 = n4920 | n4922 ;
  assign n4924 = n523 & n2558 ;
  assign n6631 = ~n4924 ;
  assign n4925 = n1052 & n6631 ;
  assign n4926 = n5595 & n4924 ;
  assign n6632 = ~n4926 ;
  assign n4927 = n2567 & n6632 ;
  assign n6633 = ~n4925 ;
  assign n4928 = n6633 & n4927 ;
  assign n6634 = ~n4928 ;
  assign n4929 = n2567 & n6634 ;
  assign n4930 = n4926 | n4928 ;
  assign n4931 = n4925 | n4930 ;
  assign n6635 = ~n4929 ;
  assign n4932 = n6635 & n4931 ;
  assign n6636 = ~n4923 ;
  assign n4933 = n6636 & n4932 ;
  assign n6637 = ~n4932 ;
  assign n4934 = n4923 & n6637 ;
  assign n4935 = n4933 | n4934 ;
  assign n3382 = n2713 & n6278 ;
  assign n3342 = n2831 & n3335 ;
  assign n3348 = n2693 & n6272 ;
  assign n4936 = n3342 | n3348 ;
  assign n4937 = n2699 & n3314 ;
  assign n4938 = n4936 | n4937 ;
  assign n4939 = n3382 | n4938 ;
  assign n6638 = ~n4939 ;
  assign n4940 = n523 & n6638 ;
  assign n4941 = n5542 & n4939 ;
  assign n4942 = n4940 | n4941 ;
  assign n6639 = ~n4942 ;
  assign n4943 = n4935 & n6639 ;
  assign n6640 = ~n4935 ;
  assign n4944 = n6640 & n4942 ;
  assign n4945 = n4943 | n4944 ;
  assign n4946 = n4860 & n4867 ;
  assign n6641 = ~n4946 ;
  assign n4947 = n4859 & n6641 ;
  assign n3949 = n2748 & n6409 ;
  assign n4948 = n2733 & n3673 ;
  assign n4949 = n2742 & n6372 ;
  assign n4950 = n4948 | n4949 ;
  assign n4951 = n3949 | n4950 ;
  assign n4952 = n2727 & n3965 ;
  assign n4953 = n4951 | n4952 ;
  assign n4954 = n672 & n4953 ;
  assign n4955 = n672 | n4953 ;
  assign n6642 = ~n4954 ;
  assign n4956 = n6642 & n4955 ;
  assign n4958 = n4947 | n4956 ;
  assign n4959 = n4947 & n4956 ;
  assign n6643 = ~n4959 ;
  assign n4960 = n4958 & n6643 ;
  assign n4961 = n4945 | n4960 ;
  assign n4962 = n4945 & n6643 ;
  assign n4963 = n4958 & n4962 ;
  assign n6644 = ~n4963 ;
  assign n4964 = n4961 & n6644 ;
  assign n4965 = n4919 & n4964 ;
  assign n4966 = n4919 | n4964 ;
  assign n6645 = ~n4965 ;
  assign n4967 = n6645 & n4966 ;
  assign n4968 = n4917 & n4967 ;
  assign n4969 = n4917 | n4967 ;
  assign n6646 = ~n4968 ;
  assign n4970 = n6646 & n4969 ;
  assign n6647 = ~n4915 ;
  assign n4971 = n6647 & n4970 ;
  assign n6648 = ~n4970 ;
  assign n4972 = n4915 & n6648 ;
  assign n4973 = n4971 | n4972 ;
  assign n4974 = n4904 | n4973 ;
  assign n4975 = n4904 & n4973 ;
  assign n6649 = ~n4975 ;
  assign n4976 = n4974 & n6649 ;
  assign n4977 = n4895 & n4976 ;
  assign n4978 = n4895 | n4976 ;
  assign n6650 = ~n4977 ;
  assign n4979 = n6650 & n4978 ;
  assign n4980 = n4897 | n4898 ;
  assign n4981 = n4077 & n4980 ;
  assign n4982 = n4979 & n4981 ;
  assign n4983 = n4979 | n4981 ;
  assign n6651 = ~n4982 ;
  assign n35 = n6651 & n4983 ;
  assign n4985 = n4915 & n4970 ;
  assign n4986 = n4975 | n4985 ;
  assign n4987 = n937 | n995 ;
  assign n4988 = n498 | n4987 ;
  assign n4989 = n3791 | n4988 ;
  assign n4990 = n635 | n4989 ;
  assign n4991 = n452 | n4990 ;
  assign n4992 = n333 | n4991 ;
  assign n4993 = n4965 | n4968 ;
  assign n6652 = ~n4947 ;
  assign n4957 = n6652 & n4956 ;
  assign n6653 = ~n4957 ;
  assign n4994 = n6653 & n4961 ;
  assign n4119 = n2727 & n4115 ;
  assign n5015 = n2733 & n6372 ;
  assign n5016 = n2742 & n6409 ;
  assign n5017 = n5015 | n5016 ;
  assign n5018 = n4119 | n5017 ;
  assign n5019 = n672 | n5018 ;
  assign n5020 = n672 & n5018 ;
  assign n6654 = ~n5020 ;
  assign n5021 = n5019 & n6654 ;
  assign n4995 = n4934 | n4944 ;
  assign n4996 = n523 & n3335 ;
  assign n6655 = ~n4930 ;
  assign n4997 = n6655 & n4996 ;
  assign n6656 = ~n4996 ;
  assign n4998 = n4930 & n6656 ;
  assign n4999 = n4997 | n4998 ;
  assign n3681 = n2699 & n3673 ;
  assign n5000 = n2693 & n3314 ;
  assign n5001 = n2831 & n6272 ;
  assign n5002 = n5000 | n5001 ;
  assign n5003 = n3681 | n5002 ;
  assign n5004 = n2713 & n3696 ;
  assign n5005 = n5003 | n5004 ;
  assign n5006 = n523 & n5005 ;
  assign n5007 = n523 | n5005 ;
  assign n6657 = ~n5006 ;
  assign n5008 = n6657 & n5007 ;
  assign n5009 = n4999 & n5008 ;
  assign n5011 = n4999 | n5008 ;
  assign n6658 = ~n5009 ;
  assign n5012 = n6658 & n5011 ;
  assign n5013 = n4995 | n5012 ;
  assign n5014 = n4995 & n5012 ;
  assign n6659 = ~n5014 ;
  assign n5022 = n5013 & n6659 ;
  assign n6660 = ~n5022 ;
  assign n5023 = n5021 & n6660 ;
  assign n6661 = ~n5021 ;
  assign n5024 = n5013 & n6661 ;
  assign n5025 = n6659 & n5024 ;
  assign n5026 = n5023 | n5025 ;
  assign n5027 = n4994 & n5026 ;
  assign n5028 = n4994 | n5026 ;
  assign n6662 = ~n5027 ;
  assign n5029 = n6662 & n5028 ;
  assign n6663 = ~n4993 ;
  assign n5030 = n6663 & n5029 ;
  assign n6664 = ~n5029 ;
  assign n5031 = n4993 & n6664 ;
  assign n5032 = n5030 | n5031 ;
  assign n5033 = n4992 & n5032 ;
  assign n5034 = n4992 | n5032 ;
  assign n6665 = ~n5033 ;
  assign n5035 = n6665 & n5034 ;
  assign n6666 = ~n4986 ;
  assign n5036 = n6666 & n5035 ;
  assign n6667 = ~n5035 ;
  assign n5037 = n4986 & n6667 ;
  assign n5038 = n5036 | n5037 ;
  assign n5039 = n4977 & n5038 ;
  assign n5040 = n4977 | n5038 ;
  assign n6668 = ~n5039 ;
  assign n5041 = n6668 & n5040 ;
  assign n5042 = n4979 | n4980 ;
  assign n5043 = n4077 & n5042 ;
  assign n5044 = n5041 & n5043 ;
  assign n5045 = n5041 | n5043 ;
  assign n6669 = ~n5044 ;
  assign n36 = n6669 & n5045 ;
  assign n5047 = n4986 & n5035 ;
  assign n5048 = n5033 | n5047 ;
  assign n5049 = n174 | n183 ;
  assign n5050 = n205 | n5049 ;
  assign n5051 = n232 | n5050 ;
  assign n5052 = n332 | n5051 ;
  assign n5053 = n2371 | n5052 ;
  assign n5054 = n972 | n5053 ;
  assign n5055 = n4087 | n5054 ;
  assign n5056 = n2252 | n5055 ;
  assign n5057 = n377 | n5056 ;
  assign n5058 = n136 | n5057 ;
  assign n5059 = n131 | n5058 ;
  assign n5060 = n209 | n5059 ;
  assign n5061 = n4993 & n5029 ;
  assign n6670 = ~n5061 ;
  assign n5062 = n5028 & n6670 ;
  assign n6671 = ~n5012 ;
  assign n5063 = n4995 & n6671 ;
  assign n5064 = n5023 | n5063 ;
  assign n3954 = n2733 & n6409 ;
  assign n4113 = n2727 & n6468 ;
  assign n5065 = n3954 | n4113 ;
  assign n6672 = ~n5065 ;
  assign n5066 = n672 & n6672 ;
  assign n5067 = n5514 & n5065 ;
  assign n5068 = n5066 | n5067 ;
  assign n3828 = n2713 & n6375 ;
  assign n3320 = n2831 & n3314 ;
  assign n3682 = n2693 & n3673 ;
  assign n5069 = n3320 | n3682 ;
  assign n5070 = n2699 & n6372 ;
  assign n5071 = n5069 | n5070 ;
  assign n5072 = n3828 | n5071 ;
  assign n6673 = ~n5072 ;
  assign n5073 = n523 & n6673 ;
  assign n5074 = n5542 & n5072 ;
  assign n5075 = n5073 | n5074 ;
  assign n6674 = ~n5075 ;
  assign n5076 = n5068 & n6674 ;
  assign n6675 = ~n5068 ;
  assign n5077 = n6675 & n5075 ;
  assign n5078 = n5076 | n5077 ;
  assign n5079 = n523 & n6272 ;
  assign n6676 = ~n5079 ;
  assign n5080 = n4996 & n6676 ;
  assign n5082 = n6656 & n5079 ;
  assign n5083 = n5080 | n5082 ;
  assign n6677 = ~n4999 ;
  assign n5010 = n6677 & n5008 ;
  assign n5084 = n4998 | n5010 ;
  assign n5085 = n5083 & n5084 ;
  assign n6678 = ~n5082 ;
  assign n5086 = n6678 & n5084 ;
  assign n5087 = n5080 | n5086 ;
  assign n5088 = n5082 | n5087 ;
  assign n6679 = ~n5085 ;
  assign n5089 = n6679 & n5088 ;
  assign n5090 = n5078 & n5089 ;
  assign n5091 = n5078 | n5089 ;
  assign n6680 = ~n5090 ;
  assign n5092 = n6680 & n5091 ;
  assign n6681 = ~n5064 ;
  assign n5093 = n6681 & n5092 ;
  assign n6682 = ~n5092 ;
  assign n5094 = n5064 & n6682 ;
  assign n5095 = n5093 | n5094 ;
  assign n5096 = n5062 | n5095 ;
  assign n5097 = n5062 & n5095 ;
  assign n6683 = ~n5097 ;
  assign n5098 = n5096 & n6683 ;
  assign n6684 = ~n5060 ;
  assign n5099 = n6684 & n5098 ;
  assign n6685 = ~n5098 ;
  assign n5100 = n5060 & n6685 ;
  assign n5101 = n5099 | n5100 ;
  assign n6686 = ~n5101 ;
  assign n5102 = n5048 & n6686 ;
  assign n6687 = ~n5048 ;
  assign n5103 = n6687 & n5101 ;
  assign n5104 = n5102 | n5103 ;
  assign n5105 = n5039 & n5104 ;
  assign n5106 = n5039 | n5104 ;
  assign n6688 = ~n5105 ;
  assign n5107 = n6688 & n5106 ;
  assign n5108 = n5041 | n5042 ;
  assign n5109 = n4077 & n5108 ;
  assign n5110 = n5107 & n5109 ;
  assign n5111 = n5107 | n5109 ;
  assign n6689 = ~n5110 ;
  assign n37 = n6689 & n5111 ;
  assign n5113 = n5060 & n5098 ;
  assign n5114 = n5048 & n5101 ;
  assign n5115 = n5113 | n5114 ;
  assign n5116 = n192 | n391 ;
  assign n5117 = n253 | n5116 ;
  assign n5118 = n357 | n5117 ;
  assign n5119 = n114 | n5118 ;
  assign n5120 = n153 | n5119 ;
  assign n5121 = n4053 | n5120 ;
  assign n5122 = n308 | n5121 ;
  assign n5123 = n2179 | n5122 ;
  assign n5124 = n1006 | n5123 ;
  assign n5125 = n3758 | n5124 ;
  assign n5126 = n194 | n5125 ;
  assign n5127 = n340 | n5126 ;
  assign n5128 = n255 | n5127 ;
  assign n5129 = n166 | n5128 ;
  assign n5130 = n139 | n5129 ;
  assign n5131 = n469 | n5130 ;
  assign n5132 = n348 | n5131 ;
  assign n6690 = ~n5094 ;
  assign n5133 = n6690 & n5096 ;
  assign n3968 = n2713 & n3965 ;
  assign n3683 = n2831 & n3673 ;
  assign n3812 = n2693 & n6372 ;
  assign n5134 = n3683 | n3812 ;
  assign n5135 = n2699 & n6409 ;
  assign n5136 = n5134 | n5135 ;
  assign n5137 = n3968 | n5136 ;
  assign n6691 = ~n5137 ;
  assign n5138 = n523 & n6691 ;
  assign n5139 = n5542 & n5137 ;
  assign n5140 = n5138 | n5139 ;
  assign n3322 = n523 & n3314 ;
  assign n5081 = n672 & n6676 ;
  assign n5141 = n5514 & n5079 ;
  assign n5142 = n5081 | n5141 ;
  assign n6692 = ~n5142 ;
  assign n5143 = n3322 & n6692 ;
  assign n6693 = ~n3322 ;
  assign n5144 = n6693 & n5142 ;
  assign n5145 = n5143 | n5144 ;
  assign n5146 = n5140 | n5145 ;
  assign n5147 = n5140 & n5145 ;
  assign n6694 = ~n5147 ;
  assign n5148 = n5146 & n6694 ;
  assign n6695 = ~n5087 ;
  assign n5149 = n6695 & n5148 ;
  assign n6696 = ~n5148 ;
  assign n5150 = n5087 & n6696 ;
  assign n5151 = n5149 | n5150 ;
  assign n5152 = n5068 & n5075 ;
  assign n6697 = ~n5089 ;
  assign n5153 = n5078 & n6697 ;
  assign n5154 = n5152 | n5153 ;
  assign n6698 = ~n5154 ;
  assign n5155 = n5151 & n6698 ;
  assign n6699 = ~n5151 ;
  assign n5156 = n6699 & n5154 ;
  assign n5157 = n5155 | n5156 ;
  assign n6700 = ~n5157 ;
  assign n5158 = n5133 & n6700 ;
  assign n6701 = ~n5133 ;
  assign n5159 = n6701 & n5157 ;
  assign n5160 = n5158 | n5159 ;
  assign n5162 = n5132 & n5160 ;
  assign n5161 = n5132 | n5160 ;
  assign n5163 = n5115 & n5161 ;
  assign n6702 = ~n5162 ;
  assign n5164 = n6702 & n5163 ;
  assign n6703 = ~n5164 ;
  assign n5165 = n5115 & n6703 ;
  assign n5166 = n5162 | n5163 ;
  assign n6704 = ~n5166 ;
  assign n5167 = n5161 & n6704 ;
  assign n5168 = n5165 | n5167 ;
  assign n5169 = n5105 | n5168 ;
  assign n5170 = n5105 & n5168 ;
  assign n6705 = ~n5170 ;
  assign n5171 = n5169 & n6705 ;
  assign n5172 = n5107 | n5108 ;
  assign n5173 = n4077 & n5172 ;
  assign n5174 = n5171 & n5173 ;
  assign n5175 = n5171 | n5173 ;
  assign n6706 = ~n5174 ;
  assign n38 = n6706 & n5175 ;
  assign n5177 = n2371 | n2438 ;
  assign n5178 = n472 | n5177 ;
  assign n5179 = n993 | n5178 ;
  assign n5180 = n2191 | n5179 ;
  assign n5181 = n1514 | n5180 ;
  assign n5182 = n1009 | n5181 ;
  assign n5183 = n3301 | n5182 ;
  assign n5184 = n135 | n5183 ;
  assign n5185 = n173 | n5184 ;
  assign n5186 = n124 | n5185 ;
  assign n5187 = n340 | n5186 ;
  assign n5188 = n367 | n5187 ;
  assign n5189 = n333 | n5188 ;
  assign n5190 = n505 | n5189 ;
  assign n5191 = n4556 & n4620 ;
  assign n5192 = n4619 | n5191 ;
  assign n5193 = n4699 & n5192 ;
  assign n5194 = n4698 | n5193 ;
  assign n5195 = n4809 & n5194 ;
  assign n5196 = n4808 | n5195 ;
  assign n5197 = n4884 & n5196 ;
  assign n5198 = n4883 | n5197 ;
  assign n5199 = n4966 & n5198 ;
  assign n5200 = n4965 | n5199 ;
  assign n5201 = n5029 & n5200 ;
  assign n6707 = ~n5201 ;
  assign n5202 = n5028 & n6707 ;
  assign n5203 = n5095 | n5202 ;
  assign n5204 = n6690 & n5203 ;
  assign n5205 = n5157 | n5204 ;
  assign n6708 = ~n5156 ;
  assign n5206 = n6708 & n5205 ;
  assign n6709 = ~n5145 ;
  assign n5207 = n5140 & n6709 ;
  assign n5208 = n5150 | n5207 ;
  assign n5209 = n523 & n3673 ;
  assign n5211 = n5141 | n5143 ;
  assign n6710 = ~n5211 ;
  assign n5212 = n5209 & n6710 ;
  assign n6711 = ~n5209 ;
  assign n5213 = n6711 & n5211 ;
  assign n5214 = n5212 | n5213 ;
  assign n3813 = n2831 & n6372 ;
  assign n3955 = n2693 & n6409 ;
  assign n5215 = n3813 | n3955 ;
  assign n5216 = n2713 & n4115 ;
  assign n5217 = n5215 | n5216 ;
  assign n5218 = n523 & n5217 ;
  assign n5219 = n523 | n5217 ;
  assign n6712 = ~n5218 ;
  assign n5220 = n6712 & n5219 ;
  assign n6713 = ~n5214 ;
  assign n5221 = n6713 & n5220 ;
  assign n6714 = ~n5220 ;
  assign n5222 = n5214 & n6714 ;
  assign n5223 = n5221 | n5222 ;
  assign n6715 = ~n5223 ;
  assign n5224 = n5208 & n6715 ;
  assign n6716 = ~n5208 ;
  assign n5225 = n6716 & n5223 ;
  assign n5226 = n5224 | n5225 ;
  assign n6717 = ~n5226 ;
  assign n5227 = n5206 & n6717 ;
  assign n6718 = ~n5206 ;
  assign n5228 = n6718 & n5226 ;
  assign n5229 = n5227 | n5228 ;
  assign n6719 = ~n5190 ;
  assign n5230 = n6719 & n5229 ;
  assign n6720 = ~n5229 ;
  assign n5231 = n5190 & n6720 ;
  assign n5232 = n5230 | n5231 ;
  assign n5233 = n5166 | n5232 ;
  assign n5234 = n5166 & n5232 ;
  assign n6721 = ~n5234 ;
  assign n5235 = n5233 & n6721 ;
  assign n5236 = n5170 & n5235 ;
  assign n5237 = n5170 | n5235 ;
  assign n6722 = ~n5236 ;
  assign n5238 = n6722 & n5237 ;
  assign n5239 = n5171 | n5172 ;
  assign n5240 = n4077 & n5239 ;
  assign n5241 = n5238 & n5240 ;
  assign n5242 = n5238 | n5240 ;
  assign n6723 = ~n5241 ;
  assign n39 = n6723 & n5242 ;
  assign n5244 = n5190 & n5229 ;
  assign n5245 = n5234 | n5244 ;
  assign n5246 = n334 | n1193 ;
  assign n5247 = n325 | n5246 ;
  assign n5248 = n252 | n5247 ;
  assign n5249 = n996 | n5248 ;
  assign n5250 = n341 | n5249 ;
  assign n5251 = n5052 | n5250 ;
  assign n5252 = n2379 | n5251 ;
  assign n5253 = n1162 | n5252 ;
  assign n5254 = n124 | n5253 ;
  assign n5255 = n224 | n5254 ;
  assign n5256 = n215 | n5255 ;
  assign n5257 = n353 | n5256 ;
  assign n5258 = n505 | n5257 ;
  assign n5259 = n752 | n5258 ;
  assign n3956 = n2831 & n6409 ;
  assign n4114 = n2713 & n6468 ;
  assign n5260 = n3956 | n4114 ;
  assign n6724 = ~n5260 ;
  assign n5261 = n523 & n6724 ;
  assign n5262 = n5542 & n5260 ;
  assign n5263 = n5261 | n5262 ;
  assign n5264 = n523 & n6374 ;
  assign n5265 = n5263 & n5264 ;
  assign n5266 = n5263 | n5264 ;
  assign n6725 = ~n5265 ;
  assign n5267 = n6725 & n5266 ;
  assign n5268 = n5213 | n5221 ;
  assign n6726 = ~n5268 ;
  assign n5269 = n5267 & n6726 ;
  assign n6727 = ~n5267 ;
  assign n5270 = n6727 & n5268 ;
  assign n5271 = n5269 | n5270 ;
  assign n5272 = n5133 | n5157 ;
  assign n5273 = n6708 & n5272 ;
  assign n5274 = n5226 | n5273 ;
  assign n6728 = ~n5224 ;
  assign n5275 = n6728 & n5274 ;
  assign n5276 = n5271 & n5275 ;
  assign n5277 = n5271 | n5275 ;
  assign n6729 = ~n5276 ;
  assign n5278 = n6729 & n5277 ;
  assign n5280 = n5259 & n5278 ;
  assign n5279 = n5259 | n5278 ;
  assign n5281 = n5245 & n5279 ;
  assign n6730 = ~n5280 ;
  assign n5282 = n6730 & n5281 ;
  assign n6731 = ~n5282 ;
  assign n5283 = n5245 & n6731 ;
  assign n5284 = n5280 | n5281 ;
  assign n6732 = ~n5284 ;
  assign n5285 = n5279 & n6732 ;
  assign n5286 = n5283 | n5285 ;
  assign n5287 = n5236 | n5286 ;
  assign n5288 = n5236 & n5286 ;
  assign n6733 = ~n5288 ;
  assign n5289 = n5287 & n6733 ;
  assign n5290 = n5238 | n5239 ;
  assign n5291 = n4077 & n5290 ;
  assign n5292 = n5289 & n5291 ;
  assign n5293 = n5289 | n5291 ;
  assign n6734 = ~n5292 ;
  assign n40 = n6734 & n5293 ;
  assign n5295 = n637 | n2316 ;
  assign n5296 = n2254 | n5295 ;
  assign n5297 = n5119 | n5296 ;
  assign n5298 = n231 | n5297 ;
  assign n5299 = n474 | n5298 ;
  assign n5300 = n3761 | n5299 ;
  assign n5301 = n206 | n5300 ;
  assign n5302 = n446 | n5301 ;
  assign n5303 = n476 | n5302 ;
  assign n6735 = ~n5270 ;
  assign n5304 = n6735 & n5277 ;
  assign n6736 = ~n5264 ;
  assign n5305 = n5263 & n6736 ;
  assign n5306 = n3807 | n5209 ;
  assign n6737 = ~n5306 ;
  assign n5307 = n523 & n6737 ;
  assign n5308 = n5305 | n5307 ;
  assign n5309 = n5304 | n5308 ;
  assign n5310 = n5304 & n5308 ;
  assign n6738 = ~n5310 ;
  assign n5311 = n5309 & n6738 ;
  assign n5210 = n6409 & n5209 ;
  assign n5312 = n3947 & n6711 ;
  assign n5313 = n5210 | n5312 ;
  assign n5314 = n523 & n5313 ;
  assign n6739 = ~n5311 ;
  assign n5315 = n6739 & n5314 ;
  assign n6740 = ~n5314 ;
  assign n5316 = n5311 & n6740 ;
  assign n5317 = n5315 | n5316 ;
  assign n5318 = n5303 | n5317 ;
  assign n5319 = n5303 & n5317 ;
  assign n6741 = ~n5319 ;
  assign n5320 = n5318 & n6741 ;
  assign n6742 = ~n5320 ;
  assign n5321 = n5284 & n6742 ;
  assign n5322 = n5284 & n5318 ;
  assign n5323 = n5319 | n5322 ;
  assign n6743 = ~n5323 ;
  assign n5324 = n5318 & n6743 ;
  assign n5325 = n5321 | n5324 ;
  assign n5326 = n5288 | n5325 ;
  assign n5327 = n5288 & n5325 ;
  assign n6744 = ~n5327 ;
  assign n5328 = n5326 & n6744 ;
  assign n5329 = n5289 | n5290 ;
  assign n5330 = n4077 & n5329 ;
  assign n5331 = n5328 & n5330 ;
  assign n5332 = n5328 | n5330 ;
  assign n6745 = ~n5331 ;
  assign n41 = n6745 & n5332 ;
  assign n5334 = n155 | n791 ;
  assign n5335 = n932 | n5334 ;
  assign n5336 = n257 | n5335 ;
  assign n5337 = n3285 | n5336 ;
  assign n5338 = n570 | n5337 ;
  assign n5339 = n1006 | n5338 ;
  assign n5340 = n136 | n5339 ;
  assign n5341 = n205 | n5340 ;
  assign n5342 = n294 | n5341 ;
  assign n5343 = n365 | n5342 ;
  assign n5344 = n213 | n5343 ;
  assign n5345 = n5323 | n5344 ;
  assign n5346 = n5323 & n5344 ;
  assign n6746 = ~n5346 ;
  assign n5347 = n5345 & n6746 ;
  assign n6747 = ~n5347 ;
  assign n5348 = n5327 & n6747 ;
  assign n5349 = n6744 & n5347 ;
  assign n5350 = n5348 | n5349 ;
  assign n5351 = n5328 | n5329 ;
  assign n5352 = n4077 & n5351 ;
  assign n5353 = n5350 & n5352 ;
  assign n5354 = n5350 | n5352 ;
  assign n6748 = ~n5353 ;
  assign n42 = n6748 & n5354 ;
  assign n5356 = n5327 & n5347 ;
  assign n5357 = n587 | n2171 ;
  assign n5358 = n607 | n5357 ;
  assign n5359 = n1200 | n5358 ;
  assign n5360 = n1155 | n5359 ;
  assign n5361 = n1012 | n5360 ;
  assign n5362 = n3733 | n5361 ;
  assign n5363 = n173 | n5362 ;
  assign n5364 = n225 | n5363 ;
  assign n5365 = n205 | n5364 ;
  assign n5366 = n354 | n5365 ;
  assign n5367 = n236 | n5366 ;
  assign n5368 = n5346 | n5367 ;
  assign n6749 = ~n5368 ;
  assign n5369 = n5356 & n6749 ;
  assign n5370 = n5346 & n5367 ;
  assign n6750 = ~n5370 ;
  assign n5371 = n5368 & n6750 ;
  assign n6751 = ~n5356 ;
  assign n5372 = n6751 & n5371 ;
  assign n5373 = n5369 | n5372 ;
  assign n5374 = n5350 | n5351 ;
  assign n5375 = n4077 & n5374 ;
  assign n5376 = n5373 & n5375 ;
  assign n5377 = n5373 | n5375 ;
  assign n6752 = ~n5376 ;
  assign n43 = n6752 & n5377 ;
  assign n5379 = n5356 & n5368 ;
  assign n5380 = n4427 | n5248 ;
  assign n5381 = n370 | n5380 ;
  assign n5382 = n2544 | n5381 ;
  assign n5383 = n964 | n5382 ;
  assign n5384 = n141 | n5383 ;
  assign n5385 = n149 | n5384 ;
  assign n5386 = n206 | n5385 ;
  assign n5387 = n137 | n5386 ;
  assign n5388 = n445 | n5387 ;
  assign n5389 = n295 | n5388 ;
  assign n5390 = n204 | n5389 ;
  assign n5391 = n5370 | n5390 ;
  assign n5392 = n5370 & n5390 ;
  assign n6753 = ~n5392 ;
  assign n5393 = n5391 & n6753 ;
  assign n5394 = n5379 & n5393 ;
  assign n5395 = n5379 | n5393 ;
  assign n6754 = ~n5394 ;
  assign n5396 = n6754 & n5395 ;
  assign n5397 = n5373 | n5374 ;
  assign n5398 = n4077 & n5397 ;
  assign n5399 = n5396 & n5398 ;
  assign n5400 = n5396 | n5398 ;
  assign n6755 = ~n5399 ;
  assign n44 = n6755 & n5400 ;
  assign n5402 = n187 | n458 ;
  assign n5403 = n1025 | n5402 ;
  assign n5404 = n501 | n5403 ;
  assign n5405 = n4742 | n5404 ;
  assign n5406 = n366 | n5405 ;
  assign n5407 = n192 | n5406 ;
  assign n5408 = n225 | n5407 ;
  assign n5409 = n309 | n5408 ;
  assign n5410 = n216 | n5409 ;
  assign n5411 = n211 | n5410 ;
  assign n5412 = n210 | n5411 ;
  assign n5413 = n553 | n5412 ;
  assign n5414 = n5392 | n5413 ;
  assign n6756 = ~n5414 ;
  assign n5415 = n5394 & n6756 ;
  assign n5416 = n5392 & n5413 ;
  assign n6757 = ~n5416 ;
  assign n5417 = n5414 & n6757 ;
  assign n5418 = n6754 & n5417 ;
  assign n5419 = n5415 | n5418 ;
  assign n5420 = n5396 | n5397 ;
  assign n5421 = n4077 & n5420 ;
  assign n5422 = n5419 & n5421 ;
  assign n5423 = n5419 | n5421 ;
  assign n6758 = ~n5422 ;
  assign n45 = n6758 & n5423 ;
  assign n5425 = n5394 & n5414 ;
  assign n5426 = n488 | n3662 ;
  assign n5427 = n441 | n5426 ;
  assign n5428 = n340 | n5427 ;
  assign n5429 = n357 | n5428 ;
  assign n5430 = n5416 | n5429 ;
  assign n5431 = n5416 & n5429 ;
  assign n6759 = ~n5431 ;
  assign n5432 = n5430 & n6759 ;
  assign n6760 = ~n5425 ;
  assign n5433 = n6760 & n5432 ;
  assign n6761 = ~n5432 ;
  assign n5434 = n5425 & n6761 ;
  assign n5435 = n5433 | n5434 ;
  assign n5436 = n5419 | n5420 ;
  assign n5437 = n4077 & n5436 ;
  assign n5438 = n5435 & n5437 ;
  assign n5439 = n5435 | n5437 ;
  assign n6762 = ~n5438 ;
  assign n46 = n6762 & n5439 ;
  assign n5441 = n5425 & n5432 ;
  assign n5442 = n441 | n516 ;
  assign n5443 = n5431 | n5442 ;
  assign n5444 = n5441 & n5443 ;
  assign n5445 = n5431 & n5442 ;
  assign n6763 = ~n5445 ;
  assign n5446 = n5443 & n6763 ;
  assign n5447 = n5441 | n5446 ;
  assign n6764 = ~n5444 ;
  assign n5448 = n6764 & n5447 ;
  assign n5449 = n5435 | n5436 ;
  assign n5451 = n4077 & n5449 ;
  assign n5452 = n5448 | n5451 ;
  assign n5453 = n5448 & n5451 ;
  assign n6765 = ~n5453 ;
  assign n47 = n5452 & n6765 ;
  assign n69 = x[21] | n67 ;
  assign n5455 = x[22] | n69 ;
  assign n5456 = n6764 & n5445 ;
  assign n5457 = n5444 & n6763 ;
  assign n5458 = n5456 | n5457 ;
  assign n5450 = n5448 | n5449 ;
  assign n5459 = n4077 & n5450 ;
  assign n5460 = n5458 & n5459 ;
  assign n5461 = n5458 | n5459 ;
  assign n6766 = ~n5460 ;
  assign n5462 = n6766 & n5461 ;
  assign n6767 = ~n5462 ;
  assign n5463 = n5455 & n6767 ;
  assign n5464 = n5444 | n5445 ;
  assign n5465 = n5450 | n5464 ;
  assign n5466 = n5444 & n5445 ;
  assign n5467 = n5450 & n5466 ;
  assign n6768 = ~n5467 ;
  assign n5468 = n5465 & n6768 ;
  assign n6769 = ~n5468 ;
  assign n5469 = n5455 & n6769 ;
  assign n6770 = ~n5469 ;
  assign n49 = n4077 & n6770 ;
  assign n48 = ~n5463 ;
  assign y[0] = n25 ;
  assign y[1] = n26 ;
  assign y[2] = n27 ;
  assign y[3] = n28 ;
  assign y[4] = n29 ;
  assign y[5] = n30 ;
  assign y[6] = n31 ;
  assign y[7] = n32 ;
  assign y[8] = n33 ;
  assign y[9] = n34 ;
  assign y[10] = n35 ;
  assign y[11] = n36 ;
  assign y[12] = n37 ;
  assign y[13] = n38 ;
  assign y[14] = n39 ;
  assign y[15] = n40 ;
  assign y[16] = n41 ;
  assign y[17] = n42 ;
  assign y[18] = n43 ;
  assign y[19] = n44 ;
  assign y[20] = n45 ;
  assign y[21] = n46 ;
  assign y[22] = n47 ;
  assign y[23] = n48 ;
  assign y[24] = n49 ;
endmodule
